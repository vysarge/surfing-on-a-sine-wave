module shark_rom #(parameter WIDTH = 40,
                    parameter HEIGHT = 20,
                    parameter LOG_FRAMES = 3)
                   (input [5:0] x,
                   input [4:0] y,
                   input [2:0] s_type,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> (WIDTH * 12 - x*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        if (s_type == 1) begin //if coin collectable
            casex({frame,y}) 
                8'b00x_00000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b00x_00001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_000_000;
				8'b00x_00010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_acc_688_000;
				8'b00x_00011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_244_acc_acc_acc_000;
				8'b00x_00100: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_222_244_244_244_244_244_244_000_000_000_000_222_244_222_244_244_acc_acc_acc_acc_000;
				8'b00x_00101: horiz=480'h_000_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_244_244_244_244_244_244_222_244_244_622_244_244_688_acc_acc_acc_688_000;
				8'b00x_00110: horiz=480'h_000_244_244_244_000_000_000_000_000_000_000_000_000_000_000_244_244_acc_688_244_244_244_244_244_244_244_244_244_244_244_ea8_244_688_acc_acc_e22_e22_e22_e22_000;
				8'b00x_00111: horiz=480'h_000_000_244_244_244_000_000_000_000_000_000_000_000_000_244_688_688_244_244_244_244_244_244_244_244_244_244_244_244_222_688_acc_acc_e22_e22_e22_e82_e82_e82_000;
				8'b00x_01000: horiz=480'h_000_000_688_688_244_244_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_acc_acc_e22_e82_eee_eee_eee_eee_eee_eee_000;
				8'b00x_01001: horiz=480'h_000_000_000_000_000_244_244_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_688_acc_eee_eee_eee_eee_eee_eee_622_622_eee_acc_ea8;
				8'b00x_01010: horiz=480'h_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_222_244_688_688_acc_eee_eee_222_eee_622_622_eee_622_622_622_eee_000;
				8'b00x_01011: horiz=480'h_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_688_222_688_acc_222_222_222_222_222_622_622_622_622_622_acc_eee_000;
				8'b00x_01100: horiz=480'h_000_000_000_000_244_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_688_acc_e22_e22_222_222_222_622_642_622_622_622_acc_eee_000_000;
				8'b00x_01101: horiz=480'h_000_000_000_244_244_244_688_000_000_000_688_244_244_244_244_244_244_244_244_244_244_244_222_222_244_acc_e22_eee_e22_ea8_e22_622_622_622_622_acc_eee_000_000_000;
				8'b00x_01110: horiz=480'h_000_000_000_244_244_000_000_000_000_244_244_688_688_acc_acc_688_688_688_244_244_688_244_244_688_688_688_acc_eee_eee_e22_622_e22_e22_622_e22_eee_000_000_000_000;
				8'b00x_01111: horiz=480'h_000_000_244_244_000_000_000_000_688_688_000_000_000_688_acc_acc_acc_acc_acc_688_244_244_244_688_acc_acc_acc_eee_eee_e22_eee_e22_e22_622_e22_acc_eee_000_000_000;
				8'b00x_10000: horiz=480'h_000_000_688_000_000_000_000_000_000_000_000_000_000_000_000_688_acc_acc_acc_244_244_244_688_acc_acc_acc_acc_e22_acc_eee_eee_e22_e22_e22_622_622_acc_acc_000_000;
				8'b00x_10001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_244_244_688_acc_acc_acc_acc_688_acc_e22_eee_eee_eee_eee_e22_622_ea8_acc_eee_000_000;
				8'b00x_10010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_000_000_000_000_000_688_688_688_acc_e82_e22_eee_eee_eee_eee_eee_eee_000_000_000;
				8'b00x_10011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_000_000_000_000_000_000_000_000_000_000_000_688_622_e82_e82_e22_e22_e22_000_000_000_000;



				8'b01x_00000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00100: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00101: horiz=480'h_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00110: horiz=480'h_000_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00111: horiz=480'h_000_000_244_244_000_000_000_000_000_000_000_000_000_000_244_244_acc_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000;
				8'b01x_01000: horiz=480'h_000_000_244_244_244_000_000_000_000_244_000_000_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_244_688_244_000_000_000;
				8'b01x_01001: horiz=480'h_000_000_000_000_688_244_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_222_688_222_244_244_244_244_000;
				8'b01x_01010: horiz=480'h_000_000_000_244_244_244_244_244_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_222_ea8_e82_244_244_244_244_244_688;
				8'b01x_01011: horiz=480'h_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_222_244_222_244_244_acc_acc_688_244_244_688_688_acc_acc_acc_688;
				8'b01x_01100: horiz=480'h_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_222_244_688_acc_688_688_688_acc_acc_acc_acc_acc_acc_688_000;
				8'b01x_01101: horiz=480'h_000_000_000_244_244_244_244_688_000_688_244_244_244_244_244_244_244_244_244_244_244_244_244_222_244_244_acc_688_acc_eee_eee_ea8_e22_688_688_688_688_eee_eee_000;
				8'b01x_01110: horiz=480'h_000_000_000_244_244_688_000_000_000_000_244_244_688_688_244_244_244_244_244_244_244_244_244_244_222_acc_eee_e22_e22_e22_eee_e22_e22_eee_eee_acc_acc_000_000_000;
				8'b01x_01111: horiz=480'h_000_000_000_244_688_000_000_000_000_244_688_000_000_acc_acc_acc_acc_acc_acc_688_244_244_244_244_acc_acc_eee_eee_e22_e22_acc_e22_eee_000_000_000_000_000_000_000;
				8'b01x_10000: horiz=480'h_000_000_244_688_000_000_000_000_000_000_000_000_000_000_688_acc_acc_acc_acc_244_244_244_244_688_acc_acc_acc_eee_eee_e22_e22_e22_eee_eee_000_000_000_000_000_000;
				8'b01x_10001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_acc_688_244_244_244_688_acc_acc_acc_688_acc_622_eee_eee_e22_eee_000_000_000_000_000_000_000;
				8'b01x_10010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_688_688_688_688_688_acc_acc_acc_622_acc_eee_eee_000_000_000_000_000_000_000;
				8'b01x_10011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_000_000_000_000_000_000_000_000_000_688_688_acc_acc_688_000_000_000_000_000_000_000;


				8'b1xx_00000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00100: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00101: horiz=480'h_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_222_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00110: horiz=480'h_000_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00111: horiz=480'h_000_000_244_244_000_000_000_000_000_000_000_000_000_000_244_244_acc_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000;
				8'b1xx_01000: horiz=480'h_000_000_244_244_244_000_000_000_000_244_000_000_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000;
				8'b1xx_01001: horiz=480'h_000_000_000_000_688_244_244_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000;
				8'b1xx_01010: horiz=480'h_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_222_244_244_000_000_000_000;
				8'b1xx_01011: horiz=480'h_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_688_244_222_244_244_222_688_688_244_688_000_000_000;
				8'b1xx_01100: horiz=480'h_000_000_000_000_244_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_688_244_244_688_244_ea8_e82_222_244_244_244_000;
				8'b1xx_01101: horiz=480'h_000_000_000_244_244_688_000_000_000_000_244_244_688_688_244_244_244_244_244_244_244_244_244_244_244_244_244_222_244_688_acc_eee_eee_acc_acc_688_688_688_acc_688;
				8'b1xx_01110: horiz=480'h_000_000_000_244_688_000_000_000_000_244_688_000_000_acc_acc_acc_acc_acc_acc_688_244_244_244_244_244_244_688_688_688_acc_acc_acc_ec4_eee_eee_acc_acc_688_688_000;
				8'b1xx_01111: horiz=480'h_000_000_244_688_000_000_000_000_000_000_000_000_000_000_688_acc_acc_acc_acc_244_244_244_244_244_244_acc_acc_acc_acc_acc_acc_acc_acc_acc_acc_000_000_000_000_000;
				8'b1xx_10000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_688_688_244_244_244_244_688_acc_acc_acc_acc_acc_688_688_acc_acc_000_000_000_000_000_000_000;
				8'b1xx_10001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_acc_acc_acc_acc_acc_acc_acc_688_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_10010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_10011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;

                
                default: horiz = 480'h_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        end
        else begin
            horiz = 0;
        end
    end
    
endmodule

module heart_rom #(parameter WIDTH = 80,
                    parameter HEIGHT = 80,
                    parameter LOG_FRAMES = 1)
                   (input [10:0] x,
                   input [9:0] y,
                   input [2:0] s_type,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> ((WIDTH  - (x>>3))*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        casex({frame,y[6:3]}) 
        	5'b0_0000: horiz=120'h_000_222_222_222_000_000_222_222_222_000;
			5'b0_0001: horiz=120'h_222_733_a23_b23_222_322_a23_b23_633_222;
			5'b0_0010: horiz=120'h_122_923_b22_b22_221_311_b22_b22_823_122;
			5'b0_0011: horiz=120'h_122_923_b22_b22_b22_b22_b22_b22_823_122;
			5'b0_0100: horiz=120'h_122_923_b22_b22_b22_b22_b22_b22_823_212;
			5'b0_0101: horiz=120'h_121_823_923_b22_b22_b22_b22_933_623_211;
			5'b0_0110: horiz=120'h_000_222_221_c12_b22_c12_c12_221_222_000;
			5'b0_0111: horiz=120'h_000_000_000_212_b23_a23_122_000_000_000;
			5'b0_1000: horiz=120'h_000_000_000_ccc_411_412_ccc_000_000_000;
			5'b0_1001: horiz=120'h_000_000_000_000_211_222_000_000_000_000;

			5'b1_0000: horiz=120'h_000_112_222_222_000_000_222_222_555_000;
			5'b1_0001: horiz=120'h_222_ccc_ccc_bbb_222_222_ccc_ccc_666_222;
			5'b1_0010: horiz=120'h_222_999_000_000_222_222_000_000_999_222;
			5'b1_0011: horiz=120'h_222_000_000_000_000_000_000_000_999_222;
			5'b1_0100: horiz=120'h_222_000_000_000_000_000_000_000_999_222;
			5'b1_0101: horiz=120'h_222_000_000_000_000_000_000_000_999_222;
			5'b1_0110: horiz=120'h_000_222_222_000_000_000_000_222_555_000;
			5'b1_0111: horiz=120'h_000_000_000_222_000_000_222_000_000_000;
			5'b1_1000: horiz=120'h_000_000_000_222_000_000_222_000_000_000;
			5'b1_1001: horiz=120'h_000_000_000_000_222_222_000_000_000_000;

			default: horiz=0;
		endcase
	end
endmodule

module number_rom #(parameter WIDTH = 40,
                    parameter HEIGHT = 50,
                    parameter LOG_FRAMES = 4)
                   (input [10:0] x,
                   input [9:0] y,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[(WIDTH>>2)*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> ((WIDTH  - (x>>2))*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        casex({frame,y[5:2]}) 
        	9'b0000_0000: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0000_0001: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0000_0010: horiz=108'h_000_111_111_000_000_000_111_111_111;
			9'b0000_0011: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_0100: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_0101: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_0110: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_0111: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_1000: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_1001: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_1010: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0000_1011: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0000_1100: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0001_0000: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_0001: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_0010: horiz=108'h_000_000_000_000_000_111_111_111_000;
			9'b0001_0011: horiz=108'h_000_000_000_111_111_111_111_111_000;
			9'b0001_0100: horiz=108'h_000_000_000_111_111_000_111_111_000;
			9'b0001_0101: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_0110: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_0111: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_1000: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_1001: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_1010: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_1011: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0001_1100: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0010_0000: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0010_0001: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0010_0010: horiz=108'h_000_111_111_000_000_000_111_111_111;
			9'b0010_0011: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0010_0100: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0010_0101: horiz=108'h_000_000_000_000_000_111_111_000_000;
			9'b0010_0110: horiz=108'h_000_000_000_000_111_111_111_000_000;
			9'b0010_0111: horiz=108'h_000_000_000_000_111_000_000_000_000;
			9'b0010_1000: horiz=108'h_000_000_111_111_000_000_000_000_000;
			9'b0010_1001: horiz=108'h_000_111_111_111_000_000_000_000_000;
			9'b0010_1010: horiz=108'h_000_111_000_000_000_000_000_000_000;
			9'b0010_1011: horiz=108'h_000_111_111_111_111_111_111_111_111;
			9'b0010_1100: horiz=108'h_000_111_111_111_111_111_111_111_000;
			9'b0011_0000: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0011_0001: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0011_0010: horiz=108'h_000_111_111_000_000_000_111_111_111;
			9'b0011_0011: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0011_0100: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0011_0101: horiz=108'h_000_000_000_000_111_111_111_000_000;
			9'b0011_0110: horiz=108'h_000_000_000_000_111_111_111_111_000;
			9'b0011_0111: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0011_1000: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0011_1001: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b0011_1010: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b0011_1011: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0011_1100: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0100_0000: horiz=108'h_000_000_000_000_000_000_111_000_000;
			9'b0100_0001: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0100_0010: horiz=108'h_000_000_000_000_111_111_111_111_000;
			9'b0100_0011: horiz=108'h_000_000_000_111_111_111_111_111_000;
			9'b0100_0100: horiz=108'h_000_000_000_111_111_000_111_111_000;
			9'b0100_0101: horiz=108'h_000_111_111_000_000_000_111_111_000;
			9'b0100_0110: horiz=108'h_111_111_111_000_000_000_111_111_000;
			9'b0100_0111: horiz=108'h_111_000_000_000_000_000_111_000_000;
			9'b0100_1000: horiz=108'h_111_111_111_111_111_111_111_111_111;
			9'b0100_1001: horiz=108'h_111_111_111_111_111_111_111_111_111;
			9'b0100_1010: horiz=108'h_000_000_000_000_000_000_111_000_000;
			9'b0100_1011: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0100_1100: horiz=108'h_000_000_000_000_000_000_111_111_000;
			9'b0101_0000: horiz=108'h_000_111_111_111_111_111_111_111_000;
			9'b0101_0001: horiz=108'h_000_111_111_111_111_111_111_111_111;
			9'b0101_0010: horiz=108'h_000_111_111_000_000_000_000_000_000;
			9'b0101_0011: horiz=108'h_000_111_111_000_000_000_000_000_000;
			9'b0101_0100: horiz=108'h_000_111_000_000_000_000_000_000_000;
			9'b0101_0101: horiz=108'h_000_111_111_111_111_111_111_000_000;
			9'b0101_0110: horiz=108'h_000_111_111_111_111_111_111_111_000;
			9'b0101_0111: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0101_1000: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0101_1001: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b0101_1010: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b0101_1011: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0101_1100: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0110_0000: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0110_0001: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0110_0010: horiz=108'h_000_111_111_000_000_000_111_111_111;
			9'b0110_0011: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0110_0100: horiz=108'h_000_111_111_000_000_000_000_000_000;
			9'b0110_0101: horiz=108'h_000_111_111_000_111_111_111_000_000;
			9'b0110_0110: horiz=108'h_000_111_111_111_111_111_111_111_000;
			9'b0110_0111: horiz=108'h_000_111_111_111_000_000_000_111_111;
			9'b0110_1000: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0110_1001: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b0110_1010: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b0110_1011: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0110_1100: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b0111_0000: horiz=108'h_000_111_111_111_111_111_111_111_000;
			9'b0111_0001: horiz=108'h_000_111_111_111_111_111_111_111_111;
			9'b0111_0010: horiz=108'h_000_000_000_000_000_000_111_111_111;
			9'b0111_0011: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0111_0100: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b0111_0101: horiz=108'h_000_000_000_000_000_111_111_000_000;
			9'b0111_0110: horiz=108'h_000_000_000_000_000_111_111_000_000;
			9'b0111_0111: horiz=108'h_000_000_000_000_000_111_111_000_000;
			9'b0111_1000: horiz=108'h_000_000_000_000_111_111_000_000_000;
			9'b0111_1001: horiz=108'h_000_000_000_000_111_111_000_000_000;
			9'b0111_1010: horiz=108'h_000_000_000_000_111_111_000_000_000;
			9'b0111_1011: horiz=108'h_000_000_000_000_111_111_000_000_000;
			9'b0111_1100: horiz=108'h_000_000_000_000_111_111_000_000_000;
			9'b1000_0000: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1000_0001: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1000_0010: horiz=108'h_000_111_111_000_000_000_111_111_111;
			9'b1000_0011: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b1000_0100: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b1000_0101: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1000_0110: horiz=108'h_000_111_111_111_111_111_111_111_000;
			9'b1000_0111: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b1000_1000: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b1000_1001: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b1000_1010: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b1000_1011: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1000_1100: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1001_0000: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1001_0001: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1001_0010: horiz=108'h_000_111_111_000_000_000_111_111_111;
			9'b1001_0011: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b1001_0100: horiz=108'h_000_111_111_000_000_000_000_111_111;
			9'b1001_0101: horiz=108'h_000_111_111_000_000_111_111_111_111;
			9'b1001_0110: horiz=108'h_000_111_111_111_111_111_111_111_111;
			9'b1001_0111: horiz=108'h_000_000_111_111_111_000_000_111_111;
			9'b1001_1000: horiz=108'h_000_000_000_000_000_000_000_111_111;
			9'b1001_1001: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b1001_1010: horiz=108'h_000_111_000_000_000_000_000_111_111;
			9'b1001_1011: horiz=108'h_000_000_111_111_111_111_111_000_000;
			9'b1001_1100: horiz=108'h_000_000_111_111_111_111_111_000_000;

			default: horiz=108'h_F00_F00_F00_F00_F00_F00_F00_F00_F00;
		endcase
	end
endmodule