`timescale 1ns / 1ps


////////////////////////////////////////////////////////////////////////////
//
//  Module that will output 12-bit RGB for a given x and y and frame and sprite type
//  Values hard-coded below.
//  s_type = 0, collectable
//           4, character
//
////////////////////////////////////////////////////////////////////////////
module sprite_rom #(parameter WIDTH = 20,
                    parameter HEIGHT = 20,
                    parameter LOG_FRAMES = 3)
                   (input [4:0] x, //height and width are both 20
                   input [4:0] y,
                   input [2:0] s_type,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> (WIDTH * 12 - x*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    /*always @(x, horiz) begin
        case (x) 
            5'b00000: pixel = horiz[239:228];
            5'b00001: pixel = horiz[227:216];
            5'b00010: pixel = horiz[215:204];
            5'b00011: pixel = horiz[203:192];
            5'b00100: pixel = horiz[191:180];
            5'b00101: pixel = horiz[179:168];
            5'b00110: pixel = horiz[167:156];
            5'b00111: pixel = horiz[155:144];
            5'b01000: pixel = horiz[143:132];
            5'b01001: pixel = horiz[131:120];
            5'b01010: pixel = horiz[119:108];
            5'b01011: pixel = horiz[107:96];
            5'b01100: pixel = horiz[95:84];
            5'b01101: pixel = horiz[83:72];
            5'b01110: pixel = horiz[71:60];
            5'b01111: pixel = horiz[59:48];
            5'b10000: pixel = horiz[47:36];
            5'b10001: pixel = horiz[35:24];
            5'b10010: pixel = horiz[23:12];
            5'b10011: pixel = horiz[11:0];
        endcase
    end*/
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        
        
        ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
        // 20 wide, 20 tall
        //
        if (s_type == 3'b100) begin //character sprite
            case ({frame,y})
                8'b000_00000: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00001: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00010: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00011: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00100: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00101: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00110: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_00111: horiz = 240'h000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000;
                8'b000_01000: horiz = 240'h000_000_0F0_0F0_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000;
                8'b000_01001: horiz = 240'h000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000;
                8'b000_01010: horiz = 240'h000_000_0F0_0F0_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000;
                8'b000_01011: horiz = 240'h000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000;
                8'b000_01100: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_01101: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_01110: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_01111: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_10000: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_10001: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_10010: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b000_10011: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                
                8'b001_00000: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_00001: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_00010: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_00011: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b001_00100: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b001_00101: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b001_00110: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b001_00111: horiz = 240'h000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000;
                8'b001_01000: horiz = 240'h000_000_0F0_0F0_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000;
                8'b001_01001: horiz = 240'h000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000;
                8'b001_01010: horiz = 240'h000_000_0F0_0F0_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000;
                8'b001_01011: horiz = 240'h000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000;
                8'b001_01100: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b001_01101: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_01110: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_01111: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_10000: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_10001: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_10010: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b001_10011: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                
                8'b010_00000: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00001: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00010: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00011: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00100: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00101: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00110: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_00111: horiz = 240'h000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000;
                8'b010_01000: horiz = 240'h000_000_0F0_0F0_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000;
                8'b010_01001: horiz = 240'h000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000;
                8'b010_01010: horiz = 240'h000_000_0F0_0F0_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000;
                8'b010_01011: horiz = 240'h000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000;
                8'b010_01100: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b010_01101: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b010_01110: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b010_01111: horiz = 240'h000_000_000_000_000_000_000_0F0_0F0_0F0_0F0_0F0_0F0_000_000_000_000_000_000_000;
                8'b010_10000: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_10001: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_10010: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b010_10011: horiz = 240'h000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                
                
                default: horiz = 240'hF00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        end
        
        
        
        //////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
        //  15 wide, 16 tall
        else if (s_type == 0) begin //collectable sprite
            case({frame,y})
                8'b000_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b000_00001: horiz = 180'h000_000_000_111_111_B70_D92_EC2_D92_B70_111_111_000_000_000;
                8'b000_00010: horiz = 180'h000_000_111_B70_EC2_EC2_EC2_EC2_EC2_EC2_EC2_B70_111_000_000;
                8'b000_00011: horiz = 180'h000_111_B70_EC2_EC2_D92_D92_D92_D92_EC2_EC2_EC2_B70_111_000;
                8'b000_00100: horiz = 180'h000_111_EC2_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_EC2_111_000;
                8'b000_00101: horiz = 180'h111_B70_EC2_D92_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_B70_111;
                8'b000_00110: horiz = 180'h111_D92_EC2_D92_D92_EC2_D92_EC2_D92_EC2_D92_FD3_EC2_D92_111;
                8'b000_00111: horiz = 180'h111_D92_EC2_D92_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_D92_111;
                8'b000_01000: horiz = 180'h111_D92_EC2_D92_D92_EC2_D92_EC2_D92_EC2_D92_FD3_EC2_D92_111;
                8'b000_01001: horiz = 180'h111_D92_EC2_D92_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_D92_111;
                8'b000_01010: horiz = 180'h111_B70_EC2_EC2_D92_EC2_D92_EC2_D92_EC2_EC2_FD3_EC2_B70_111;
                8'b000_01011: horiz = 180'h000_111_EC2_EC2_FD3_D92_EC2_D92_EC2_EC2_FD3_EC2_EC2_111_000;
                8'b000_01100: horiz = 180'h000_111_B70_EC2_EC2_FD3_FD3_FD3_FD3_FD3_EC2_EC2_B70_111_000;
                8'b000_01101: horiz = 180'h000_000_111_B70_EC2_EC2_EC2_EC2_EC2_EC2_EC2_B70_111_000_000;
                8'b000_01110: horiz = 180'h000_000_000_111_111_B70_D92_EC2_D92_B70_111_111_000_000_000;
                8'b000_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                
                8'b001_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b001_00001: horiz = 180'h000_000_000_111_111_FF4_EC2_D92_B70_950_111_111_000_000_000;
                8'b001_00010: horiz = 180'h000_000_111_D92_FFF_EC2_D92_D92_D92_D92_B70_950_111_000_000;
                8'b001_00011: horiz = 180'h000_111_D92_FFF_EC2_D92_D92_B70_B70_D92_D92_D92_950_111_000;
                8'b001_00100: horiz = 180'h000_111_FFF_FF4_D92_D92_B70_D92_B70_D92_EC2_D92_D92_111_000;
                8'b001_00101: horiz = 180'h111_D92_FF4_EC2_D92_B70_D92_B70_D92_B70_D92_EC2_D92_950_111;
                8'b001_00110: horiz = 180'h111_FF4_FF4_EC2_D92_B70_B70_D92_B70_D92_B70_EC2_D92_B70_111;
                8'b001_00111: horiz = 180'h111_ED3_ED3_D92_D92_B70_D92_B70_D92_B70_D92_EC2_D92_B70_111;
                8'b001_01000: horiz = 180'h111_EC2_EC2_D92_D92_B70_B70_D92_B70_D92_B70_EC2_D92_B70_111;
                8'b001_01001: horiz = 180'h111_D92_D92_D92_D92_B70_D92_B70_D92_B70_D92_EC2_D92_B70_111;
                8'b001_01010: horiz = 180'h111_D92_EC2_EC2_D92_D92_B70_D92_B70_D92_B70_EC2_D92_950_111;
                8'b001_01011: horiz = 180'h000_111_ED3_ED3_D92_D92_EC2_D92_D92_B70_EC2_D92_B70_111_000;
                8'b001_01100: horiz = 180'h000_111_D92_FF4_EC2_D92_D92_EC2_EC2_EC2_D92_D92_950_111_000;
                8'b001_01101: horiz = 180'h000_000_111_D92_ED3_EC2_D92_D92_D92_D92_B70_950_111_000_000;
                8'b001_01110: horiz = 180'h000_000_000_111_111_EC2_EC2_D92_B70_950_111_111_000_000_000;
                8'b001_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b010_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b010_00001: horiz = 180'h000_000_000_000_111_D92_ED3_D92_B70_740_111_000_000_000_000;
                8'b010_00010: horiz = 180'h000_000_000_111_ED3_FFF_D92_B70_B70_B70_950_111_000_000_000;
                8'b010_00011: horiz = 180'h000_000_111_D92_FFF_D92_B70_950_B70_B70_B70_740_111_000_000;
                8'b010_00100: horiz = 180'h000_000_111_ED3_FF4_B70_950_B70_950_D92_B70_950_111_000_000;
                8'b010_00101: horiz = 180'h000_111_D92_FF4_D92_B70_950_950_B70_B70_D92_B70_740_111_000;
                8'b010_00110: horiz = 180'h000_111_ED3_ED3_D92_B70_950_B70_950_B70_D92_B70_950_111_000;
                8'b010_00111: horiz = 180'h000_111_EC2_EC2_B70_B70_950_950_B70_950_D92_B70_950_111_000;
                8'b010_01000: horiz = 180'h000_111_D92_D92_B70_B70_950_B70_950_B70_D92_B70_950_111_000;
                8'b010_01001: horiz = 180'h000_111_B70_B70_B70_B70_950_950_B70_950_D92_B70_950_111_000;
                8'b010_01010: horiz = 180'h000_111_D92_D92_D92_B70_B70_B70_950_B70_D92_B70_740_111_000;
                8'b010_01011: horiz = 180'h000_000_111_EC2_EC2_B70_D92_950_B70_D92_B70_950_111_000_000;
                8'b010_01100: horiz = 180'h000_000_111_D92_ED3_D92_B70_D92_D92_B70_B70_740_111_000_000;
                8'b010_01101: horiz = 180'h000_000_000_111_EC2_EC2_D92_B70_B70_B70_950_111_000_000_000;
                8'b010_01110: horiz = 180'h000_000_000_000_111_D92_D92_D92_B70_740_111_000_000_000_000;
                8'b010_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b011_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b011_00001: horiz = 180'h000_000_000_000_111_B70_EC2_D92_B70_950_111_000_000_000_000;
                8'b011_00010: horiz = 180'h000_000_000_111_B70_ED3_ED3_B70_950_950_740_111_000_000_000;
                8'b011_00011: horiz = 180'h000_000_000_111_FF4_FFF_EC2_950_950_740_950_111_000_000_000;
                8'b011_00100: horiz = 180'h000_000_111_B70_FF4_FF4_D92_950_740_950_950_740_111_000_000;
                8'b011_00101: horiz = 180'h000_000_111_EC2_ED3_ED3_B70_950_740_740_B70_950_111_000_000;
                8'b011_00110: horiz = 180'h000_000_111_EC2_EC2_EC2_950_950_740_950_B70_950_111_000_000;
                8'b011_00111: horiz = 180'h000_000_111_D92_D92_D92_950_950_740_740_B70_950_111_000_000;
                8'b011_01000: horiz = 180'h000_000_111_B70_B70_B70_950_950_740_950_B70_950_111_000_000;
                8'b011_01001: horiz = 180'h000_000_111_950_950_950_950_950_740_740_B70_950_111_000_000;
                8'b011_01010: horiz = 180'h000_000_111_B70_B70_B70_B70_950_740_950_B70_950_111_000_000;
                8'b011_01011: horiz = 180'h000_000_111_B70_D92_D92_D92_950_950_950_B70_740_111_000_000;
                8'b011_01100: horiz = 180'h000_000_000_111_EC2_EC2_EC2_950_950_B70_950_111_000_000_000;
                8'b011_01101: horiz = 180'h000_000_000_111_B70_D92_D92_B70_950_950_740_111_000_000_000;
                8'b011_01110: horiz = 180'h000_000_000_000_111_B70_B70_D92_B70_950_111_000_000_000_000;
                8'b011_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b100_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b100_00001: horiz = 180'h000_000_000_000_000_111_EC2_EC2_EC2_111_000_000_000_000_000;
                8'b100_00010: horiz = 180'h000_000_000_000_000_111_ED3_ED3_ED3_111_000_000_000_000_000;
                8'b100_00011: horiz = 180'h000_000_000_000_000_111_FF4_FF4_FF4_111_000_000_000_000_000;
                8'b100_00100: horiz = 180'h000_000_000_000_000_111_ED3_ED3_ED3_111_000_000_000_000_000;
                8'b100_00101: horiz = 180'h000_000_000_000_000_111_EC2_EC2_EC2_111_000_000_000_000_000;
                8'b100_00110: horiz = 180'h000_000_000_000_000_111_E92_E92_E92_111_000_000_000_000_000;
                8'b100_00111: horiz = 180'h000_000_000_000_000_111_B70_B70_B70_111_000_000_000_000_000;
                8'b100_01000: horiz = 180'h000_000_000_000_000_111_950_950_950_111_000_000_000_000_000;
                8'b100_01001: horiz = 180'h000_000_000_000_000_111_740_740_740_111_000_000_000_000_000;
                8'b100_01010: horiz = 180'h000_000_000_000_000_111_950_950_950_111_000_000_000_000_000;
                8'b100_01011: horiz = 180'h000_000_000_000_000_111_B70_B70_B70_111_000_000_000_000_000;
                8'b100_01100: horiz = 180'h000_000_000_000_000_111_E92_E92_E92_111_000_000_000_000_000;
                8'b100_01101: horiz = 180'h000_000_000_000_000_111_B70_B70_B70_111_000_000_000_000_000;
                8'b100_01110: horiz = 180'h000_000_000_000_000_111_950_950_950_111_000_000_000_000_000;
                8'b100_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                

                8'b101_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b101_00001: horiz = 180'h000_000_000_000_111_EC2_ED3_D92_D92_950_111_000_000_000_000;
                8'b101_00010: horiz = 180'h000_000_000_111_EC2_FF4_FF4_ED3_EC2_EC2_740_111_000_000_000;
                8'b101_00011: horiz = 180'h000_000_000_111_ED3_FF4_FF4_FF4_ED3_ED3_D92_111_000_000_000;
                8'b101_00100: horiz = 180'h000_000_111_D92_FF4_ED3_ED3_FF4_ED3_EC2_EC2_740_111_000_000;
                8'b101_00101: horiz = 180'h000_000_111_EC2_FF4_ED3_FF4_FFF_FF4_D92_D92_950_111_000_000;
                8'b101_00110: horiz = 180'h000_000_111_ED3_FF4_ED3_ED3_FFF_FF4_B70_B70_B70_111_000_000;
                8'b101_00111: horiz = 180'h000_000_111_ED3_FF4_ED3_FF4_FFF_FF4_950_950_950_111_000_000;
                8'b101_01000: horiz = 180'h000_000_111_ED3_FF4_ED3_ED3_FFF_FF4_740_740_740_111_000_000;
                8'b101_01001: horiz = 180'h000_000_111_ED3_FF4_ED3_FF4_FFF_FF4_740_740_740_111_000_000;
                8'b101_01010: horiz = 180'h000_000_111_EC2_FF4_ED3_FF4_FFF_EC2_740_740_740_111_000_000;
                8'b101_01011: horiz = 180'h000_000_111_D92_FF4_FF4_FFF_FF4_D92_950_950_740_111_000_000;
                8'b101_01100: horiz = 180'h000_000_000_111_ED3_FF4_FF4_FF4_B70_B70_B70_111_000_000_000;
                8'b101_01101: horiz = 180'h000_000_000_111_EC2_FF4_FF4_EC2_950_950_740_111_000_000_000;
                8'b101_01110: horiz = 180'h000_000_000_000_111_EC2_FF4_D92_740_740_111_000_000_000_000;
                8'b101_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b110_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b110_00001: horiz = 180'h000_000_000_000_111_D92_FF4_ED3_D92_950_111_000_000_000_000;
                8'b110_00010: horiz = 180'h000_000_000_111_EC2_FF4_FF4_FF4_FF4_D92_950_111_000_000_000;
                8'b110_00011: horiz = 180'h000_000_111_D92_FF4_ED3_FF4_FF4_FF4_ED3_B70_740_111_000_000;
                8'b110_00100: horiz = 180'h000_000_111_ED3_ED3_FF4_ED3_FFF_FF4_FF4_D92_950_111_000_000;
                8'b110_00101: horiz = 180'h000_111_D92_FF4_ED3_ED3_FF4_FF4_FFF_FF4_EC2_D92_740_111_000;
                8'b110_00110: horiz = 180'h000_111_EC2_FF4_ED3_FF4_ED3_FF4_FFF_FF4_FF4_B70_B70_111_000;
                8'b110_00111: horiz = 180'h000_111_ED3_FF4_ED3_ED3_FF4_ED3_FFF_FF4_FF4_950_950_111_000;
                8'b110_01000: horiz = 180'h000_111_ED3_FF4_ED3_FF4_ED3_FF4_FFF_FF4_FF4_740_740_111_000;
                8'b110_01001: horiz = 180'h000_111_EC2_FF4_ED3_ED3_FF4_ED3_FFF_FF4_FF4_740_740_111_000;
                8'b110_01010: horiz = 180'h000_111_D92_FF4_ED3_FF4_ED3_FF4_FFF_FF4_EC2_740_740_111_000;
                8'b110_01011: horiz = 180'h000_000_111_ED3_FF4_ED3_FF4_FFF_FF4_FF4_D92_950_111_000_000;
                8'b110_01100: horiz = 180'h000_000_111_D92_FF4_FFF_FFF_FF4_FF4_ED3_950_740_111_000_000;
                8'b110_01101: horiz = 180'h000_000_000_111_EC2_FF4_FF4_FF4_FF4_D92_950_111_000_000_000;
                8'b110_01110: horiz = 180'h000_000_000_000_111_D92_FF4_ED3_D92_740_111_000_000_000_000;
                8'b110_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b111_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b111_00001: horiz = 180'h000_000_000_111_111_D92_ED3_ED3_D92_950_111_111_000_000_000;
                8'b111_00010: horiz = 180'h000_000_111_B70_EC2_ED3_ED3_ED3_ED3_ED3_950_740_111_000_000;
                8'b111_00011: horiz = 180'h000_111_B70_ED3_ED3_EC2_EC2_ED3_ED3_ED3_D92_D92_740_111_000;
                8'b111_00100: horiz = 180'h000_111_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_ED3_B70_B70_111_000;
                8'b111_00101: horiz = 180'h111_B70_ED3_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_D92_B70_740_111;
                8'b111_00110: horiz = 180'h111_EC2_ED3_EC2_EC2_ED3_EC2_ED3_EC2_FF4_ED3_EC2_950_950_111;
                8'b111_00111: horiz = 180'h111_EC2_ED3_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_EC2_740_740_111;
                8'b111_01000: horiz = 180'h111_EC2_ED3_EC2_EC2_ED3_EC2_ED3_EC2_FF4_ED3_EC2_740_740_111;
                8'b111_01001: horiz = 180'h111_EC2_ED3_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_EC2_740_740_111;
                8'b111_01010: horiz = 180'h111_B70_ED3_ED3_EC2_ED3_EC2_ED3_ED3_FF4_ED3_D92_740_740_111;
                8'b111_01011: horiz = 180'h000_111_EC2_ED3_FF4_ED3_ED3_ED3_FF4_ED3_ED3_950_740_111_000;
                8'b111_01100: horiz = 180'h000_111_B70_ED3_ED3_FF4_FF4_FF4_ED3_ED3_D92_740_740_111_000;
                8'b111_01101: horiz = 180'h000_000_111_B70_EC2_ED3_ED3_ED3_ED3_EC2_950_740_111_000_000;
                8'b111_01110: horiz = 180'h000_000_000_111_111_D92_ED3_ED3_D92_950_111_111_000_000_000;
                8'b111_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                
                default: horiz = 240'hF00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        end
        else begin
            horiz = 0;
        end
    end
    
endmodule

