module background_rom #(parameter WIDTH = 1024,
                    parameter HEIGHT = 512)
                   (input [10:0] x,
                   input [9:0] y,
                   output reg [11:0]  pixel);
    
    reg[(WIDTH>>4)*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = horiz >> (12*((WIDTH - x)>>4)-2);
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y, return the corresponding pixel strip
    always @(y) begin
        case(y[8:4]) 
            8'b00000: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00001: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00010: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7cf_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00011: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cd_eee_fff_eff_cef_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8ce_8cf_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00100: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6cf_7cf_7cf_7ce_7cf_7cf_7cf_7cf_abc_fff_eff_fff_fff_fff_eff_cef_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6cf_7cf_9ce_eef_fff_fff_fff_bff_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00101: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6ce_8cd_dff_efe_fff_8ce_7cf_7cf_8cd_eef_eef_eef_fff_fff_fff_fff_fff_cff_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_9ce_eef_eef_dee_fff_eff_fff_fff_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00110: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_7cf_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6cf_8ce_fff_fff_fff_fff_fff_fff_8be_def_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_eff_cff_7ce_8cf_7cf_7cf_7ce_7cf_8ce_eef_eef_eef_eef_eef_eee_fff_eff_9ce_8cd_7cf_7cf_8cf_7cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_7cf_8cf_8cf_7cf_8cf_7ce_7cf_7cf_8cf_7cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b00111: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8ce_8cd_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_def_eef_dee_fff_fff_fff_efe_def_eef_eef_eef_eef_eef_eef_fff_fff_dee_fff_fff_ffe_fff_7ce_7cf_7cf_7cf_7ce_7cf_abd_eef_eef_eee_fff_eef_eef_eef_eef_eef_eff_fff_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cd_eef_fff_eff_cef_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b01000: horiz=1536'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_6cf_8ce_9bd_eef_fff_eff_fff_cff_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_eef_eef_eef_eee_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_7ce_7ce_7cf_7cf_7cf_7cf_eef_eef_eef_eee_fff_fff_eef_eef_eee_fff_fff_fff_eff_ddf_8cd_6cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_7cf_7cf_7cf_7ce_7ce_7ce_7cf_abc_fff_eff_fff_fff_fff_eff_cef_8cf_7ce_7ce_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
			8'b01001: horiz=1536'h_7ce_7cf_7ce_7cf_7ce_7cf_7ce_7cf_7ce_7cf_7ce_7cf_7ce_7cf_7ce_7cf_7ce_7cf_7ce_8cf_7cf_9cd_eef_eef_eef_fff_eff_fff_fff_8cf_7cf_7cf_7ce_7cf_7ce_8cf_7ce_7cf_7ce_7cf_7ce_7cf_7cf_7cf_7cf_def_eef_eef_eef_eef_eef_eef_eef_eef_def_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_def_7ce_7cf_7ce_8cf_7ce_7cf_9cd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_def_eee_def_7ce_7cf_7ce_7cf_7be_7ce_9cd_def_eff_fff_9cf_7cf_7bf_9ce_eef_eef_eef_fff_fff_fff_fff_fff_dff_8cd_7cf_7cf_7ce_7cf_7cf_8cf_7ce_7cf_7ce_7cf_7cf_8cf_7ce_7cf_7ce_7cf;
			8'b01010: horiz=1536'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_9cf_eef_eef_eef_eef_eef_eee_eff_eff_ace_9ce_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9ce_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_8cf_7df_8df_8cf_8cf_8cf_8df_9ce_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_cef_8cf_8cf_8cf_8cf_8cf_8df_ace_fff_fff_fff_fff_fff_fff_9cf_def_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_eff_cff_8cf_8cf_8df_8cf_8ce_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
			8'b01011: horiz=1536'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_acd_eef_eef_eee_fff_eef_eef_eef_eef_eef_eff_eff_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9ce_def_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_eee_fff_fff_eef_eef_eef_eef_eef_cef_8df_8df_8cf_8cf_8cf_9ce_def_def_ddf_ddf_def_def_def_def_ddf_ddf_def_def_cef_8cf_8cf_8cf_8cf_8cf_8df_def_eef_dee_fff_fff_fff_eff_def_eef_eef_eef_eef_eef_eef_fff_fff_eee_fff_fff_eff_eff_8cf_8cf_8cf_8df_8df_eef_cff_9ce_8df_8df_8cf_8cf_8cf_8cf;
			8'b01100: horiz=1536'h_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8df_8df_def_def_eef_eef_fff_fff_eef_eef_eef_fff_fff_fff_fff_def_9ce_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_acd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_cef_9ce_8df_8cf_9df_def_edf_eef_cef_cef_cef_ddf_ddf_ddf_ddf_cef_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_eef_eef_eef_eee_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_8df_8cf_8df_9ce_def_eef_eef_def_cff_8ce_8cf_8cf_8cf_8cf;
			8'b01101: horiz=1536'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_9de_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_eef_eef_def_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eef_eef_eef_eef_def_def_eef_eef_cef_ace_8df_8df_8cf_8cf_8df_9df_9ce_9ce_8cf_8df_8df_8df_8cf_8cf_8df_8cf_8df_8df_8cf_8cf_8cf_8cf_8df_def_eef_eef_eef_eef_eef_eef_eef_eef_def_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_8df_8cf_8cf_9bd_cef_def_cef_8df_8df_8cf_8df_8cf_8cf;
			8'b01110: horiz=1536'h_8cf_8df_8cf_8df_8cf_8df_7de_9df_9cf_9df_9ce_8cf_8cf_8df_8cf_9df_8cf_8df_8cf_8df_9ce_9ce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_efe_eff_9ce_9df_8cf_8df_8cf_8df_8cf_8df_8cf_eef_def_def_ddf_def_def_ddf_def_eef_eef_def_def_def_def_eef_eef_def_ddf_def_ddf_ddf_def_eef_cef_cef_9de_8df_7df_9ce_abc_eef_fff_fff_fff_8df_8cf_8cf_8cf_8df_8ce_9df_8ce_8df_8cf_8df_8cf_9df_8cf_8ce_def_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_9ce_8df_8cf_8df_8cf_9df_8cf_8df_8cf_9df_8cf_8df_8cf_8df;
			8'b01111: horiz=1536'h_8cf_8cf_8cf_8cf_8cf_8cf_9ce_8ce_8cf_9ce_9cd_9ce_9df_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8ce_9de_ddf_ddf_def_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_dde_fff_cff_8ce_8ce_8cf_8cf_8cf_8cf_8cf_8cf_ace_eef_ddf_def_def_ddf_ddf_def_def_ddf_def_def_ddf_def_ddf_def_def_def_ddf_ddf_ddf_def_def_def_def_def_9de_def_eef_eef_eef_fff_fff_fff_eef_9ce_9ce_8cf_8cf_8cf_8ce_8df_8cf_8cf_8cf_8cf_8cf_8ce_9ce_def_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_eee_fff_fff_eef_eef_eef_eef_eef_cef_8df_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
			8'b10000: horiz=1536'h_8cf_8cf_8df_8cf_8ce_8cf_9ce_9bd_eef_fff_fff_fff_cff_8cf_8cf_8cf_8ce_8cf_8cf_8cf_8cf_9df_cef_ddf_def_cef_cff_def_ddf_ddf_def_def_ddf_eef_fff_fff_cff_9ce_8ce_8cf_8de_8ce_8cf_8cf_8cf_8cf_8ce_8ce_ace_cef_bef_9ce_def_def_def_cef_acd_acd_9ce_9df_dff_cef_def_cef_8ce_8ce_8cf_8cf_8cf_8cf_8cf_9cd_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_9ce_9ce_9df_9cd_dee_eef_9cd_8df_8ce_8ce_8df_acd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_dff_def_9ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
			8'b10001: horiz=1536'h_8cf_8cf_8cf_8cf_8df_acd_eef_eef_def_fff_eff_fff_fff_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9ce_9cf_8cf_9cf_8df_eef_eef_eef_fff_fff_eef_eef_eef_eef_eef_fff_eff_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_9cf_8df_8cf_9ce_9ce_9ce_8cf_8df_8cf_8cf_8cf_9cf_8cf_8cf_8cf_9cf_8cf_9de_eef_eef_eef_fff_fff_eef_eef_ddf_ddf_dee_fff_eff_8cf_acd_eef_dee_fff_fff_9ce_8ce_9df_9cf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eef_eef_eef_eef_eef_def_def_eef_eef_def_9ce_9ce_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
			8'b10010: horiz=1536'h_9df_9df_9df_9df_9de_eef_eef_eef_eef_eef_dee_fff_eff_ade_ade_adf_9df_9df_9df_9df_9df_9df_9de_9df_9df_9df_9df_ade_eef_eef_eef_fff_fff_eee_eef_eef_fff_fff_eff_fff_fff_ddf_9de_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_ade_eef_eef_eef_fff_fff_dee_eef_eee_fff_fff_eff_eff_fff_eef_eef_eef_eef_fff_eef_fff_9ce_9df_def_dde_ddf_ddf_def_ddf_ddf_def_eef_eef_def_def_ddf_eef_eef_eef_def_ddf_def_ddf_def_def_eef_cef_cef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df;
			8'b10011: horiz=1536'h_9df_9df_9df_9df_acd_eef_eef_eee_fff_eef_eef_eef_eef_eef_fff_eff_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_eef_eef_eef_eef_eef_fff_eef_eef_eef_eef_dee_fff_fff_eef_eef_cff_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9de_9df_9df_9df_9df_9df_9df_9df_9df_adf_def_eef_eef_eef_eef_eee_fff_eef_eef_eef_eef_eee_fff_fff_eef_eef_eef_eef_eef_eef_eef_def_bef_ade_def_ddf_def_ddf_ddf_ddf_ddf_def_ddf_def_ddf_cdf_def_ddf_ddf_ddf_def_def_def_ddf_cef_cef_cef_ddf_cef_adf_9df_9df_9df_9df_9df_9df_9df_9df;
			8'b10100: horiz=1536'h_9df_adf_9df_9df_eef_eef_eef_eef_fff_fff_eef_eef_eee_fff_fff_fff_fff_def_ade_9df_ade_bce_dee_def_9cf_adf_9df_9df_adf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_dee_ace_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_def_eef_edf_eef_cff_9df_9df_9df_9df_adf_bde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_adf_cef_ade_cef_cef_9df_9df_9df_9df_9df_9df_bde_cdf_bef_adf_cef_def_cef_def_bde_bce_ade_9df_cef_cef_cef_cef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
			8'b10101: horiz=1536'h_9df_9df_9df_acd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_eef_eef_def_eef_eef_fff_fff_def_9df_9df_9df_9df_def_ddf_def_ddf_ddf_def_ddf_ddf_ddf_ddf_def_def_eef_dee_fff_fff_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_bde_cef_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
			8'b10110: horiz=1536'h_9de_9df_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dff_bce_eef_eef_eef_fff_eef_eef_cef_adf_adf_adf_ddf_ddf_cef_cef_cef_cdf_ddf_ddf_def_def_eef_eef_eef_eef_fff_eef_fff_ade_9ce_9df_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_ade_ddf_def_def_eef_cef_ddf_ddf_def_edf_ddf_cef_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_adf_adf_9df_adf_9df_adf_9de_adf_9de_adf_9df_9df_adf_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf;
			8'b10111: horiz=1536'h_9df_9df_ade_cef_def_def_ddf_def_ddf_ddf_ddf_ddf_def_def_ddf_def_ddf_def_cef_adf_eef_eef_eef_eef_eef_def_eee_def_adf_adf_ade_ace_9df_9df_9df_9de_ade_ace_ade_9cf_bce_eef_eef_eef_eef_eef_eef_eef_cef_ace_9ce_9de_9de_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9de_9de_adf_cef_def_cef_cef_9df_ade_9de_ade_9de_adf_9df_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9de_9df_9de_9df_9df_9de_9ce_9de_9cf_adf_bcd_def_ade_ade_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de_9df_9de;
			8'b11000: horiz=1536'h_9df_9de_9df_9de_adf_9df_ddf_ddf_def_def_ddf_def_ddf_def_def_ddf_bef_ade_9df_9df_ade_def_cef_ade_def_def_eef_eef_def_eef_bde_9de_9df_9df_9df_9df_9df_9df_9df_9de_adf_ade_bdf_9de_def_cef_eef_eef_eef_eef_def_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_bce_adf_adf_9de_9de_ade_ddf_eef_eef_def_eef_bde_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
			8'b11001: horiz=1536'h_adf_9df_adf_9df_adf_9df_ace_cef_def_bce_bdf_9de_ade_ade_ade_ade_9df_9df_adf_adf_9df_9df_9df_9df_9df_ade_def_cef_def_9de_adf_9df_adf_9df_adf_9df_adf_9df_adf_adf_ade_9df_adf_9df_9df_9de_ace_def_def_cef_ade_9de_adf_adf_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9de_def_eef_eef_def_cff_adf_9df_ade_def_cef_def_9de_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df_adf_9df;
			8'b11010: horiz=1536'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
			8'b11011: horiz=1536'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
			8'b11100: horiz=1536'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
			8'b11101: horiz=1536'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
			8'b11110: horiz=1536'h_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_adf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef_adf_bdf_bef_bef;
			8'b11111: horiz=1536'h_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade_adf_adf_ade_ade;

            
            default: horiz = 768'h_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
        endcase

    end
    
endmodule

