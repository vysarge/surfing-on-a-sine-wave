module shark_rom #(parameter WIDTH = 40,
                    parameter HEIGHT = 20,
                    parameter LOG_FRAMES = 3)
                   (input [5:0] x,
                   input [4:0] y,
                   input [2:0] s_type,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> (WIDTH * 12 - x*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        if (s_type == 1) begin //if coin collectable
            casex({frame,y}) 
                8'b00x_00000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b00x_00001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_000_000;
				8'b00x_00010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_acc_688_000;
				8'b00x_00011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_244_acc_acc_acc_000;
				8'b00x_00100: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_222_244_244_244_244_244_244_000_000_000_000_222_244_222_244_244_acc_acc_acc_acc_000;
				8'b00x_00101: horiz=480'h_000_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_244_244_244_244_244_244_222_244_244_622_244_244_688_acc_acc_acc_688_000;
				8'b00x_00110: horiz=480'h_000_244_244_244_000_000_000_000_000_000_000_000_000_000_000_244_244_acc_688_244_244_244_244_244_244_244_244_244_244_244_ea8_244_688_acc_acc_e22_e22_e22_e22_000;
				8'b00x_00111: horiz=480'h_000_000_244_244_244_000_000_000_000_000_000_000_000_000_244_688_688_244_244_244_244_244_244_244_244_244_244_244_244_222_688_acc_acc_e22_e22_e22_e82_e82_e82_000;
				8'b00x_01000: horiz=480'h_000_000_688_688_244_244_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_acc_acc_e22_e82_eee_eee_eee_eee_eee_eee_000;
				8'b00x_01001: horiz=480'h_000_000_000_000_000_244_244_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_688_acc_eee_eee_eee_eee_eee_eee_622_622_eee_acc_ea8;
				8'b00x_01010: horiz=480'h_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_222_244_688_688_acc_eee_eee_222_eee_622_622_eee_622_622_622_eee_000;
				8'b00x_01011: horiz=480'h_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_688_222_688_acc_222_222_222_222_222_622_622_622_622_622_acc_eee_000;
				8'b00x_01100: horiz=480'h_000_000_000_000_244_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_688_acc_e22_e22_222_222_222_622_642_622_622_622_acc_eee_000_000;
				8'b00x_01101: horiz=480'h_000_000_000_244_244_244_688_000_000_000_688_244_244_244_244_244_244_244_244_244_244_244_222_222_244_acc_e22_eee_e22_ea8_e22_622_622_622_622_acc_eee_000_000_000;
				8'b00x_01110: horiz=480'h_000_000_000_244_244_000_000_000_000_244_244_688_688_acc_acc_688_688_688_244_244_688_244_244_688_688_688_acc_eee_eee_e22_622_e22_e22_622_e22_eee_000_000_000_000;
				8'b00x_01111: horiz=480'h_000_000_244_244_000_000_000_000_688_688_000_000_000_688_acc_acc_acc_acc_acc_688_244_244_244_688_acc_acc_acc_eee_eee_e22_eee_e22_e22_622_e22_acc_eee_000_000_000;
				8'b00x_10000: horiz=480'h_000_000_688_000_000_000_000_000_000_000_000_000_000_000_000_688_acc_acc_acc_244_244_244_688_acc_acc_acc_acc_e22_acc_eee_eee_e22_e22_e22_622_622_acc_acc_000_000;
				8'b00x_10001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_244_244_688_acc_acc_acc_acc_688_acc_e22_eee_eee_eee_eee_e22_622_ea8_acc_eee_000_000;
				8'b00x_10010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_000_000_000_000_000_688_688_688_acc_e82_e22_eee_eee_eee_eee_eee_eee_000_000_000;
				8'b00x_10011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_000_000_000_000_000_000_000_000_000_000_000_688_622_e82_e82_e22_e22_e22_000_000_000_000;



				8'b01x_00000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00100: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00101: horiz=480'h_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00110: horiz=480'h_000_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000;
				8'b01x_00111: horiz=480'h_000_000_244_244_000_000_000_000_000_000_000_000_000_000_244_244_acc_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000;
				8'b01x_01000: horiz=480'h_000_000_244_244_244_000_000_000_000_244_000_000_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_244_688_244_000_000_000;
				8'b01x_01001: horiz=480'h_000_000_000_000_688_244_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_222_688_222_244_244_244_244_000;
				8'b01x_01010: horiz=480'h_000_000_000_244_244_244_244_244_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_222_ea8_e82_244_244_244_244_244_688;
				8'b01x_01011: horiz=480'h_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_222_244_222_244_244_acc_acc_688_244_244_688_688_acc_acc_acc_688;
				8'b01x_01100: horiz=480'h_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_222_244_688_acc_688_688_688_acc_acc_acc_acc_acc_acc_688_000;
				8'b01x_01101: horiz=480'h_000_000_000_244_244_244_244_688_000_688_244_244_244_244_244_244_244_244_244_244_244_244_244_222_244_244_acc_688_acc_eee_eee_ea8_e22_688_688_688_688_eee_eee_000;
				8'b01x_01110: horiz=480'h_000_000_000_244_244_688_000_000_000_000_244_244_688_688_244_244_244_244_244_244_244_244_244_244_222_acc_eee_e22_e22_e22_eee_e22_e22_eee_eee_acc_acc_000_000_000;
				8'b01x_01111: horiz=480'h_000_000_000_244_688_000_000_000_000_244_688_000_000_acc_acc_acc_acc_acc_acc_688_244_244_244_244_acc_acc_eee_eee_e22_e22_acc_e22_eee_000_000_000_000_000_000_000;
				8'b01x_10000: horiz=480'h_000_000_244_688_000_000_000_000_000_000_000_000_000_000_688_acc_acc_acc_acc_244_244_244_244_688_acc_acc_acc_eee_eee_e22_e22_e22_eee_eee_000_000_000_000_000_000;
				8'b01x_10001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_acc_688_244_244_244_688_acc_acc_acc_688_acc_622_eee_eee_e22_eee_000_000_000_000_000_000_000;
				8'b01x_10010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_688_688_688_688_688_acc_acc_acc_622_acc_eee_eee_000_000_000_000_000_000_000;
				8'b01x_10011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_000_000_000_000_000_000_000_000_000_688_688_acc_acc_688_000_000_000_000_000_000_000;


				8'b1xx_00000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00100: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00101: horiz=480'h_244_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_222_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00110: horiz=480'h_000_244_244_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_688_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_00111: horiz=480'h_000_000_244_244_000_000_000_000_000_000_000_000_000_000_244_244_acc_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000_000;
				8'b1xx_01000: horiz=480'h_000_000_244_244_244_000_000_000_000_244_000_000_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000_000_000;
				8'b1xx_01001: horiz=480'h_000_000_000_000_688_244_244_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_000_000_000_000_000;
				8'b1xx_01010: horiz=480'h_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_688_222_244_244_000_000_000_000;
				8'b1xx_01011: horiz=480'h_000_000_000_000_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_688_244_222_244_244_222_688_688_244_688_000_000_000;
				8'b1xx_01100: horiz=480'h_000_000_000_000_244_244_244_244_688_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_244_222_688_244_244_688_244_ea8_e82_222_244_244_244_000;
				8'b1xx_01101: horiz=480'h_000_000_000_244_244_688_000_000_000_000_244_244_688_688_244_244_244_244_244_244_244_244_244_244_244_244_244_222_244_688_acc_eee_eee_acc_acc_688_688_688_acc_688;
				8'b1xx_01110: horiz=480'h_000_000_000_244_688_000_000_000_000_244_688_000_000_acc_acc_acc_acc_acc_acc_688_244_244_244_244_244_244_688_688_688_acc_acc_acc_ec4_eee_eee_acc_acc_688_688_000;
				8'b1xx_01111: horiz=480'h_000_000_244_688_000_000_000_000_000_000_000_000_000_000_688_acc_acc_acc_acc_244_244_244_244_244_244_acc_acc_acc_acc_acc_acc_acc_acc_acc_acc_000_000_000_000_000;
				8'b1xx_10000: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_688_688_688_244_244_244_244_688_acc_acc_acc_acc_acc_688_688_acc_acc_000_000_000_000_000_000_000;
				8'b1xx_10001: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_244_244_688_acc_acc_acc_acc_acc_acc_acc_688_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_10010: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_244_688_688_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
				8'b1xx_10011: horiz=480'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;

                
                default: horiz = 480'h_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        end
        else begin
            horiz = 0;
        end
    end
    
endmodule

