`timescale 1ns / 1ps


////////////////////////////////////////////////////////////////////////////
//
//  Module that will output 12-bit RGB for a given x and y and frame and sprite type
//  Values hard-coded below.
//  s_type = 0, collectable
//           4, character
//
////////////////////////////////////////////////////////////////////////////
module sprite_rom #(parameter WIDTH = 45,
                    parameter HEIGHT = 42,
                    parameter LOG_FRAMES = 2)
                   (input [10:0] x, //height and width are both 20
                   input [9:0] y,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> (WIDTH * 12 - x*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        
        
        ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
        // 20 wide, 20 tall
        //
        //character sprite
            casex ({frame,y})
                8'b0x_000000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_b46_b46_b46_b46_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_b46_624_624_624_624_624_624_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_000111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_b46_624_000_000_624_624_624_624_624_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001000: horiz=540'h_000_000_000_000_000_000_000_000_000_b46_624_000_fff_fff_fff_000_624_624_624_000_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001001: horiz=540'h_000_000_000_000_000_000_000_000_b46_624_624_000_fff_fff_fff_fff_000_624_fff_fff_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001010: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_000_fff_fff_fff_fff_000_624_fff_fff_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001011: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_000_fff_fff_fff_000_624_fff_fff_fff_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001100: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_000_000_624_624_624_000_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001101: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_624_624_624_624_624_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001110: horiz=540'h_000_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_000_624_624_624_b46_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_001111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010000: horiz=540'h_000_000_000_000_624_624_b46_b46_000_000_000_000_000_000_bbf_bbf_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010001: horiz=540'h_000_000_000_000_624_624_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_624_624_624_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_f40_fff_fff_f40_f40_fff_fff_fff_f40_000_000_000_624_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010011: horiz=540'h_000_000_000_000_000_000_000_000_b00_b00_bbf_bbf_bbf_b00_b00_b00_bbf_bbf_b00_f40_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010100: horiz=540'h_000_000_000_000_000_000_000_000_b00_b00_bbf_bbf_bbf_b00_b00_b00_bbf_bbf_b00_b00_bbf_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010101: horiz=540'h_000_000_000_000_000_000_000_000_bbf_b00_b00_000_000_000_000_000_000_000_b00_b00_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_602_602_000_bbf_bbf_bbf_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_010111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_011000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_011001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_fff_fff_fff_fff_000;
                8'b0x_011010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_d6b_000_000_000_000_000_000_000_fd9_fd9_fd9_fd9_fd9_f40_f40_f40_f40_f40_fff_000;
                8'b0x_011011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_b46_b46_000_000_000_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000;
                8'b0x_011100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000;
                8'b0x_011101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_f40_000_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000;
                8'b0x_011110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_f40_f40_f40_b00_b00_000_000_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000;
                8'b0x_011111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_b46_b46_d6b_000_000_000_f40_f40_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_000_000_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100000: horiz=540'h_000_000_000_000_000_000_000_000_b46_624_624_624_000_000_fd9_f40_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_000_000_000_b00_b00_b00_b00_b00_b00_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100010: horiz=540'h_000_000_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100011: horiz=540'h_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100100: horiz=540'h_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100101: horiz=540'h_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100110: horiz=540'h_000_000_fd9_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_100111: horiz=540'h_000_000_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b0x_101000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                
                8'b10_000000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_b46_b46_b46_b46_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_000111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_b46_624_624_624_624_624_624_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_b46_624_624_624_624_624_624_624_624_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001001: horiz=540'h_000_000_000_000_000_000_000_000_000_624_624_624_fff_fff_fff_000_624_624_624_fff_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001010: horiz=540'h_000_000_000_000_000_000_000_000_b46_624_624_000_fff_fff_fff_fff_000_624_fff_fff_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001011: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_000_fff_fff_fff_fff_000_624_fff_fff_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001100: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_000_fff_000_624_fff_000_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001101: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_624_624_624_624_624_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001110: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_624_624_624_624_624_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_001111: horiz=540'h_000_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_000_624_624_624_b46_000_000_000_b46_b46_624_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_b46_624_624_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_bbf_bbf_000_000_000_000_000_000_000_000_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_f40_fff_fff_f40_f40_fff_fff_fff_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010100: horiz=540'h_000_000_000_000_000_b46_b46_000_b00_b00_bbf_bbf_bbf_b00_b00_b00_bbf_bbf_b00_f40_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010101: horiz=540'h_000_000_000_000_000_624_624_000_b00_b00_bbf_bbf_bbf_b00_b00_b00_bbf_bbf_b00_b00_bbf_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010110: horiz=540'h_000_000_000_000_000_000_000_000_bbf_b00_b00_000_000_000_000_000_000_000_b00_b00_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_010111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_602_602_000_bbf_bbf_bbf_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_011000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_011001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_fff_fff_fff_fff_000;
                8'b10_011010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_d6b_000_000_000_000_000_000_000_fd9_fd9_fd9_fd9_fd9_f40_f40_f40_f40_f40_fff_000;
                8'b10_011011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_b46_b46_000_000_000_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000;
                8'b10_011100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000;
                8'b10_011101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_f40_000_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000;
                8'b10_011110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_f40_f40_f40_b00_b00_000_000_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000;
                8'b10_011111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_b46_b46_d6b_000_000_000_f40_f40_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_000_000_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000;
                8'b10_100000: horiz=540'h_000_000_000_000_000_000_000_000_b46_624_624_624_000_000_fd9_f40_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_000_000_000_b00_b00_b00_b00_b00_b00_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100010: horiz=540'h_000_000_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100011: horiz=540'h_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100100: horiz=540'h_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100101: horiz=540'h_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100110: horiz=540'h_000_000_fd9_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_100111: horiz=540'h_000_000_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b10_101000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                
                8'b11_000000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_000111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_b46_b46_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_b46_b46_624_624_624_b46_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_b46_624_624_624_624_624_624_624_624_b46_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001011: horiz=540'h_000_000_000_000_000_000_000_000_000_b46_624_624_624_624_624_624_624_624_624_b46_b46_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001100: horiz=540'h_000_000_000_000_000_000_000_000_000_624_624_624_fff_fff_fff_000_624_624_624_fff_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001101: horiz=540'h_000_000_000_000_000_000_000_000_b46_624_624_000_fff_fff_fff_fff_000_624_fff_fff_000_000_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001110: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_000_fff_000_624_fff_000_b46_624_624_d6b_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_001111: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_624_624_624_624_000_624_624_624_b46_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010000: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_624_624_624_624_000_624_624_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010001: horiz=540'h_000_000_000_000_000_000_000_000_000_624_624_624_624_624_624_624_000_624_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_624_624_624_624_624_000_000_624_624_624_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_bbf_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_602_b00_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010110: horiz=540'h_000_000_000_000_000_000_000_000_000_f40_bbf_bbf_bbf_b00_b00_b00_bbf_fff_f40_f40_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_010111: horiz=540'h_000_000_000_000_000_000_000_000_b00_b00_bbf_bbf_bbf_b00_b00_b00_bbf_bbf_b00_b00_bbf_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_011000: horiz=540'h_000_000_000_000_000_000_000_000_bbf_b00_b00_bbf_bbf_b00_b00_bbf_bbf_bbf_b00_b00_bbf_fff_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_011001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_bbf_bbf_bbf_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_011010: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_011011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_fd9_fd9_fd9_fff_fff_fff_fff_000;
                8'b11_011100: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_d6b_d6b_000_000_000_000_fd9_fd9_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_000;
                8'b11_011101: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_b46_000_000_000_fd9_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000;
                8'b11_011110: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_fd9_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000;
                8'b11_011111: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_f40_f40_000_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000;
                8'b11_100000: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_d6b_d6b_000_000_000_000_f40_f40_f40_b00_b00_b00_b00_b00_000_000_000_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000;
                8'b11_100001: horiz=540'h_000_000_000_000_000_000_000_000_b46_b46_b46_624_000_000_000_f40_f40_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_000_000_000_f40_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_100010: horiz=540'h_000_000_000_000_000_000_000_000_624_624_624_000_000_fd9_fd9_000_000_000_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_b00_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_100011: horiz=540'h_000_000_000_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_b00_b00_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_100100: horiz=540'h_000_000_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_100101: horiz=540'h_000_000_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_100110: horiz=540'h_000_000_000_000_fd9_fd9_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_100111: horiz=540'h_000_000_fd9_fd9_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_101000: horiz=540'h_000_f40_f40_f40_f40_f40_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                8'b11_101001: horiz=540'h_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
                
                
                default: horiz = 540'h_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        
    end
    
endmodule

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  Module to store pixels for the collectable coin animation
//
module collectable_rom #(parameter WIDTH = 15,
                    parameter HEIGHT = 16,
                    parameter LOG_FRAMES = 3)
                   (input [4:0] x,
                   input [4:0] y,
                   input [2:0] s_type,
                   input [LOG_FRAMES-1:0] frame,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> (WIDTH * 12 - x*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        if (s_type == 0) begin //if coin collectable
            case({frame,y}) 
                8'b000_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b000_00001: horiz = 180'h000_000_000_111_111_B70_D92_EC2_D92_B70_111_111_000_000_000;
                8'b000_00010: horiz = 180'h000_000_111_B70_EC2_EC2_EC2_EC2_EC2_EC2_EC2_B70_111_000_000;
                8'b000_00011: horiz = 180'h000_111_B70_EC2_EC2_D92_D92_D92_D92_EC2_EC2_EC2_B70_111_000;
                8'b000_00100: horiz = 180'h000_111_EC2_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_EC2_111_000;
                8'b000_00101: horiz = 180'h111_B70_EC2_D92_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_B70_111;
                8'b000_00110: horiz = 180'h111_D92_EC2_D92_D92_EC2_D92_EC2_D92_EC2_D92_FD3_EC2_D92_111;
                8'b000_00111: horiz = 180'h111_D92_EC2_D92_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_D92_111;
                8'b000_01000: horiz = 180'h111_D92_EC2_D92_D92_EC2_D92_EC2_D92_EC2_D92_FD3_EC2_D92_111;
                8'b000_01001: horiz = 180'h111_D92_EC2_D92_EC2_D92_EC2_D92_EC2_D92_EC2_FD3_EC2_D92_111;
                8'b000_01010: horiz = 180'h111_B70_EC2_EC2_D92_EC2_D92_EC2_D92_EC2_EC2_FD3_EC2_B70_111;
                8'b000_01011: horiz = 180'h000_111_EC2_EC2_FD3_D92_EC2_D92_EC2_EC2_FD3_EC2_EC2_111_000;
                8'b000_01100: horiz = 180'h000_111_B70_EC2_EC2_FD3_FD3_FD3_FD3_FD3_EC2_EC2_B70_111_000;
                8'b000_01101: horiz = 180'h000_000_111_B70_EC2_EC2_EC2_EC2_EC2_EC2_EC2_B70_111_000_000;
                8'b000_01110: horiz = 180'h000_000_000_111_111_B70_D92_EC2_D92_B70_111_111_000_000_000;
                8'b000_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                
                8'b001_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b001_00001: horiz = 180'h000_000_000_111_111_FF4_EC2_D92_B70_950_111_111_000_000_000;
                8'b001_00010: horiz = 180'h000_000_111_D92_FFF_EC2_D92_D92_D92_D92_B70_950_111_000_000;
                8'b001_00011: horiz = 180'h000_111_D92_FFF_EC2_D92_D92_B70_B70_D92_D92_D92_950_111_000;
                8'b001_00100: horiz = 180'h000_111_FFF_FF4_D92_D92_B70_D92_B70_D92_EC2_D92_D92_111_000;
                8'b001_00101: horiz = 180'h111_D92_FF4_EC2_D92_B70_D92_B70_D92_B70_D92_EC2_D92_950_111;
                8'b001_00110: horiz = 180'h111_FF4_FF4_EC2_D92_B70_B70_D92_B70_D92_B70_EC2_D92_B70_111;
                8'b001_00111: horiz = 180'h111_ED3_ED3_D92_D92_B70_D92_B70_D92_B70_D92_EC2_D92_B70_111;
                8'b001_01000: horiz = 180'h111_EC2_EC2_D92_D92_B70_B70_D92_B70_D92_B70_EC2_D92_B70_111;
                8'b001_01001: horiz = 180'h111_D92_D92_D92_D92_B70_D92_B70_D92_B70_D92_EC2_D92_B70_111;
                8'b001_01010: horiz = 180'h111_D92_EC2_EC2_D92_D92_B70_D92_B70_D92_B70_EC2_D92_950_111;
                8'b001_01011: horiz = 180'h000_111_ED3_ED3_D92_D92_EC2_D92_D92_B70_EC2_D92_B70_111_000;
                8'b001_01100: horiz = 180'h000_111_D92_FF4_EC2_D92_D92_EC2_EC2_EC2_D92_D92_950_111_000;
                8'b001_01101: horiz = 180'h000_000_111_D92_ED3_EC2_D92_D92_D92_D92_B70_950_111_000_000;
                8'b001_01110: horiz = 180'h000_000_000_111_111_EC2_EC2_D92_B70_950_111_111_000_000_000;
                8'b001_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b010_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b010_00001: horiz = 180'h000_000_000_000_111_D92_ED3_D92_B70_740_111_000_000_000_000;
                8'b010_00010: horiz = 180'h000_000_000_111_ED3_FFF_D92_B70_B70_B70_950_111_000_000_000;
                8'b010_00011: horiz = 180'h000_000_111_D92_FFF_D92_B70_950_B70_B70_B70_740_111_000_000;
                8'b010_00100: horiz = 180'h000_000_111_ED3_FF4_B70_950_B70_950_D92_B70_950_111_000_000;
                8'b010_00101: horiz = 180'h000_111_D92_FF4_D92_B70_950_950_B70_B70_D92_B70_740_111_000;
                8'b010_00110: horiz = 180'h000_111_ED3_ED3_D92_B70_950_B70_950_B70_D92_B70_950_111_000;
                8'b010_00111: horiz = 180'h000_111_EC2_EC2_B70_B70_950_950_B70_950_D92_B70_950_111_000;
                8'b010_01000: horiz = 180'h000_111_D92_D92_B70_B70_950_B70_950_B70_D92_B70_950_111_000;
                8'b010_01001: horiz = 180'h000_111_B70_B70_B70_B70_950_950_B70_950_D92_B70_950_111_000;
                8'b010_01010: horiz = 180'h000_111_D92_D92_D92_B70_B70_B70_950_B70_D92_B70_740_111_000;
                8'b010_01011: horiz = 180'h000_000_111_EC2_EC2_B70_D92_950_B70_D92_B70_950_111_000_000;
                8'b010_01100: horiz = 180'h000_000_111_D92_ED3_D92_B70_D92_D92_B70_B70_740_111_000_000;
                8'b010_01101: horiz = 180'h000_000_000_111_EC2_EC2_D92_B70_B70_B70_950_111_000_000_000;
                8'b010_01110: horiz = 180'h000_000_000_000_111_D92_D92_D92_B70_740_111_000_000_000_000;
                8'b010_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b011_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b011_00001: horiz = 180'h000_000_000_000_111_B70_EC2_D92_B70_950_111_000_000_000_000;
                8'b011_00010: horiz = 180'h000_000_000_111_B70_ED3_ED3_B70_950_950_740_111_000_000_000;
                8'b011_00011: horiz = 180'h000_000_000_111_FF4_FFF_EC2_950_950_740_950_111_000_000_000;
                8'b011_00100: horiz = 180'h000_000_111_B70_FF4_FF4_D92_950_740_950_950_740_111_000_000;
                8'b011_00101: horiz = 180'h000_000_111_EC2_ED3_ED3_B70_950_740_740_B70_950_111_000_000;
                8'b011_00110: horiz = 180'h000_000_111_EC2_EC2_EC2_950_950_740_950_B70_950_111_000_000;
                8'b011_00111: horiz = 180'h000_000_111_D92_D92_D92_950_950_740_740_B70_950_111_000_000;
                8'b011_01000: horiz = 180'h000_000_111_B70_B70_B70_950_950_740_950_B70_950_111_000_000;
                8'b011_01001: horiz = 180'h000_000_111_950_950_950_950_950_740_740_B70_950_111_000_000;
                8'b011_01010: horiz = 180'h000_000_111_B70_B70_B70_B70_950_740_950_B70_950_111_000_000;
                8'b011_01011: horiz = 180'h000_000_111_B70_D92_D92_D92_950_950_950_B70_740_111_000_000;
                8'b011_01100: horiz = 180'h000_000_000_111_EC2_EC2_EC2_950_950_B70_950_111_000_000_000;
                8'b011_01101: horiz = 180'h000_000_000_111_B70_D92_D92_B70_950_950_740_111_000_000_000;
                8'b011_01110: horiz = 180'h000_000_000_000_111_B70_B70_D92_B70_950_111_000_000_000_000;
                8'b011_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b100_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b100_00001: horiz = 180'h000_000_000_000_000_111_EC2_EC2_EC2_111_000_000_000_000_000;
                8'b100_00010: horiz = 180'h000_000_000_000_000_111_ED3_ED3_ED3_111_000_000_000_000_000;
                8'b100_00011: horiz = 180'h000_000_000_000_000_111_FF4_FF4_FF4_111_000_000_000_000_000;
                8'b100_00100: horiz = 180'h000_000_000_000_000_111_ED3_ED3_ED3_111_000_000_000_000_000;
                8'b100_00101: horiz = 180'h000_000_000_000_000_111_EC2_EC2_EC2_111_000_000_000_000_000;
                8'b100_00110: horiz = 180'h000_000_000_000_000_111_E92_E92_E92_111_000_000_000_000_000;
                8'b100_00111: horiz = 180'h000_000_000_000_000_111_B70_B70_B70_111_000_000_000_000_000;
                8'b100_01000: horiz = 180'h000_000_000_000_000_111_950_950_950_111_000_000_000_000_000;
                8'b100_01001: horiz = 180'h000_000_000_000_000_111_740_740_740_111_000_000_000_000_000;
                8'b100_01010: horiz = 180'h000_000_000_000_000_111_950_950_950_111_000_000_000_000_000;
                8'b100_01011: horiz = 180'h000_000_000_000_000_111_B70_B70_B70_111_000_000_000_000_000;
                8'b100_01100: horiz = 180'h000_000_000_000_000_111_E92_E92_E92_111_000_000_000_000_000;
                8'b100_01101: horiz = 180'h000_000_000_000_000_111_B70_B70_B70_111_000_000_000_000_000;
                8'b100_01110: horiz = 180'h000_000_000_000_000_111_950_950_950_111_000_000_000_000_000;
                8'b100_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                

                8'b101_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b101_00001: horiz = 180'h000_000_000_000_111_EC2_ED3_D92_D92_950_111_000_000_000_000;
                8'b101_00010: horiz = 180'h000_000_000_111_EC2_FF4_FF4_ED3_EC2_EC2_740_111_000_000_000;
                8'b101_00011: horiz = 180'h000_000_000_111_ED3_FF4_FF4_FF4_ED3_ED3_D92_111_000_000_000;
                8'b101_00100: horiz = 180'h000_000_111_D92_FF4_ED3_ED3_FF4_ED3_EC2_EC2_740_111_000_000;
                8'b101_00101: horiz = 180'h000_000_111_EC2_FF4_ED3_FF4_FFF_FF4_D92_D92_950_111_000_000;
                8'b101_00110: horiz = 180'h000_000_111_ED3_FF4_ED3_ED3_FFF_FF4_B70_B70_B70_111_000_000;
                8'b101_00111: horiz = 180'h000_000_111_ED3_FF4_ED3_FF4_FFF_FF4_950_950_950_111_000_000;
                8'b101_01000: horiz = 180'h000_000_111_ED3_FF4_ED3_ED3_FFF_FF4_740_740_740_111_000_000;
                8'b101_01001: horiz = 180'h000_000_111_ED3_FF4_ED3_FF4_FFF_FF4_740_740_740_111_000_000;
                8'b101_01010: horiz = 180'h000_000_111_EC2_FF4_ED3_FF4_FFF_EC2_740_740_740_111_000_000;
                8'b101_01011: horiz = 180'h000_000_111_D92_FF4_FF4_FFF_FF4_D92_950_950_740_111_000_000;
                8'b101_01100: horiz = 180'h000_000_000_111_ED3_FF4_FF4_FF4_B70_B70_B70_111_000_000_000;
                8'b101_01101: horiz = 180'h000_000_000_111_EC2_FF4_FF4_EC2_950_950_740_111_000_000_000;
                8'b101_01110: horiz = 180'h000_000_000_000_111_EC2_FF4_D92_740_740_111_000_000_000_000;
                8'b101_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b110_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b110_00001: horiz = 180'h000_000_000_000_111_D92_FF4_ED3_D92_950_111_000_000_000_000;
                8'b110_00010: horiz = 180'h000_000_000_111_EC2_FF4_FF4_FF4_FF4_D92_950_111_000_000_000;
                8'b110_00011: horiz = 180'h000_000_111_D92_FF4_ED3_FF4_FF4_FF4_ED3_B70_740_111_000_000;
                8'b110_00100: horiz = 180'h000_000_111_ED3_ED3_FF4_ED3_FFF_FF4_FF4_D92_950_111_000_000;
                8'b110_00101: horiz = 180'h000_111_D92_FF4_ED3_ED3_FF4_FF4_FFF_FF4_EC2_D92_740_111_000;
                8'b110_00110: horiz = 180'h000_111_EC2_FF4_ED3_FF4_ED3_FF4_FFF_FF4_FF4_B70_B70_111_000;
                8'b110_00111: horiz = 180'h000_111_ED3_FF4_ED3_ED3_FF4_ED3_FFF_FF4_FF4_950_950_111_000;
                8'b110_01000: horiz = 180'h000_111_ED3_FF4_ED3_FF4_ED3_FF4_FFF_FF4_FF4_740_740_111_000;
                8'b110_01001: horiz = 180'h000_111_EC2_FF4_ED3_ED3_FF4_ED3_FFF_FF4_FF4_740_740_111_000;
                8'b110_01010: horiz = 180'h000_111_D92_FF4_ED3_FF4_ED3_FF4_FFF_FF4_EC2_740_740_111_000;
                8'b110_01011: horiz = 180'h000_000_111_ED3_FF4_ED3_FF4_FFF_FF4_FF4_D92_950_111_000_000;
                8'b110_01100: horiz = 180'h000_000_111_D92_FF4_FFF_FFF_FF4_FF4_ED3_950_740_111_000_000;
                8'b110_01101: horiz = 180'h000_000_000_111_EC2_FF4_FF4_FF4_FF4_D92_950_111_000_000_000;
                8'b110_01110: horiz = 180'h000_000_000_000_111_D92_FF4_ED3_D92_740_111_000_000_000_000;
                8'b110_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;

                8'b111_00000: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                8'b111_00001: horiz = 180'h000_000_000_111_111_D92_ED3_ED3_D92_950_111_111_000_000_000;
                8'b111_00010: horiz = 180'h000_000_111_B70_EC2_ED3_ED3_ED3_ED3_ED3_950_740_111_000_000;
                8'b111_00011: horiz = 180'h000_111_B70_ED3_ED3_EC2_EC2_ED3_ED3_ED3_D92_D92_740_111_000;
                8'b111_00100: horiz = 180'h000_111_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_ED3_B70_B70_111_000;
                8'b111_00101: horiz = 180'h111_B70_ED3_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_D92_B70_740_111;
                8'b111_00110: horiz = 180'h111_EC2_ED3_EC2_EC2_ED3_EC2_ED3_EC2_FF4_ED3_EC2_950_950_111;
                8'b111_00111: horiz = 180'h111_EC2_ED3_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_EC2_740_740_111;
                8'b111_01000: horiz = 180'h111_EC2_ED3_EC2_EC2_ED3_EC2_ED3_EC2_FF4_ED3_EC2_740_740_111;
                8'b111_01001: horiz = 180'h111_EC2_ED3_EC2_ED3_EC2_ED3_EC2_ED3_FF4_ED3_EC2_740_740_111;
                8'b111_01010: horiz = 180'h111_B70_ED3_ED3_EC2_ED3_EC2_ED3_ED3_FF4_ED3_D92_740_740_111;
                8'b111_01011: horiz = 180'h000_111_EC2_ED3_FF4_ED3_ED3_ED3_FF4_ED3_ED3_950_740_111_000;
                8'b111_01100: horiz = 180'h000_111_B70_ED3_ED3_FF4_FF4_FF4_ED3_ED3_D92_740_740_111_000;
                8'b111_01101: horiz = 180'h000_000_111_B70_EC2_ED3_ED3_ED3_ED3_EC2_950_740_111_000_000;
                8'b111_01110: horiz = 180'h000_000_000_111_111_D92_ED3_ED3_D92_950_111_111_000_000_000;
                8'b111_01111: horiz = 180'h000_000_000_000_000_111_111_111_111_111_000_000_000_000_000;
                
                default: horiz = 180'hF00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        end
        else begin
            horiz = 180'hFF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0;
        end
    end
    
endmodule

