module background_rom #(parameter WIDTH = 40,
                    parameter HEIGHT = 20,
                    parameter LOG_FRAMES = 3)
                   (input [10:0] x,
                   input [9:0] y,
                   input [10:0] offset,
                   output reg [11:0]  pixel);
    
    reg[WIDTH*12-1:0] horiz; //a horizontal strip of pixels
    //selects the correct pixel from the horizontal strip
    
    always @(x, horiz) begin
        pixel = (horiz >> (WIDTH * 12 - (x+offset)*12 - 12));
        //[WIDTH*12-1-x*12:WIDTH*12-13-x*12];
    end
    
    
    //for current y and frame, return the corresponding pixel strip
    always @(y, frame) begin
        if (s_type == 1) begin //if coin collectable
            case(y) 
                8'b000000000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000000111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000001111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000010111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000011111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000100111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000101111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000110111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b000111111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001000111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001001111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001010111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001011111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001100111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001101111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001110111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7df_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6cf_7cf_7cf_7cf_8df_7cf_7cf_7cf_7cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8ce_8ce_8bd_9cd_9cd_9cd_9cd_9cd_9cd_9cd_9cd_9cd_9cd_8ce_9df_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b001111111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_8ce_8ce_8cd_cff_dee_eff_eff_eff_eff_eff_eff_eff_eff_eff_eff_cff_cff_8cd_8ce_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8ce_9cd_9bc_acc_bcd_def_efe_fff_fff_fff_fff_fff_eff_eff_eff_eff_eff_dee_cee_9bc_add_8cd_8ce_8be_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7cf_7cf_7cf_7cf_7df_7cf_7cf_8ce_9ce_9cd_9cc_acc_9cc_9cd_9cc_9cd_9cd_9ce_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8ce_9de_cff_dff_eff_eff_eef_fff_fff_fff_fff_fff_fff_eff_eff_fff_eff_eff_eff_eff_eff_dff_cef_bef_8cd_8ce_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7ce_8ce_9ce_dff_dff_eff_eff_eff_eff_eff_dff_cff_cff_8bd_8cf_8cf_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8bd_9cd_9cd_dff_dee_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_eff_def_cef_9bd_9cd_9ce_8cf_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_9df_9cd_9cd_acd_def_eff_fff_eff_eff_fff_fff_eff_def_cee_9bc_9cd_9ce_8df_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000011: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_abd_dff_def_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_cff_bef_8ce_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_7cf_7ce_8ce_9ce_dff_def_def_dee_fff_fff_fff_ffe_fff_fff_fff_fff_fff_eff_fff_eff_dff_bff_7ce_7cf_7df_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000100: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7df_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8ce_9df_bcd_dff_def_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_dff_9cd_9ce_8cf_7cf_7cf_7df_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8be_8ce_8bd_9cd_8cd_9cd_bce_ddf_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_def_cff_8ce_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000101: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7df_7cf_7cf_7cf_8cf_8cf_8cf_8cf_7cf_7cf_8cf_8ce_8cf_7cf_7cf_6cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8ce_9ce_dff_def_def_eef_def_def_eef_def_dee_eee_fff_fff_eff_fff_fff_fff_fff_eff_eff_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_cff_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8cf_9ce_cef_def_cef_dff_def_eef_dde_eef_eef_dee_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_eff_eff_eff_dff_9cd_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000110: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8ce_9ce_8cd_9cd_9cd_9cd_9cd_9cd_9cd_9cd_9cd_8cd_8ce_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_9ce_acd_def_def_def_eef_ddf_eef_eef_eef_eef_eef_eff_eff_fff_fff_fff_fff_fff_fff_eff_eff_eff_eff_eff_fff_fff_eff_eff_fff_fff_fff_dff_def_ace_9cf_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7be_8ce_9ce_9ce_acd_def_dee_dde_eef_eef_eef_eef_eef_eef_dee_eff_eff_eff_eff_fff_eff_eff_eff_fff_fff_eff_fff_eff_eff_9cd_9cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010000111: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8ce_8ce_9ce_dff_dff_eff_eff_eff_eff_eff_eff_eff_eff_cef_cef_8bd_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8ce_cff_def_ede_dee_eee_eef_eef_eef_eef_eef_eef_def_dee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_ffe_fff_eff_eff_dff_cff_8ce_8ce_8cf_7cf_7cf_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7ce_8ce_cef_cef_def_def_def_eee_ede_eef_eef_eef_eef_eef_eef_eee_fff_eff_fff_fff_fff_eff_eff_fff_fff_fff_fff_fff_fff_fff_def_bef_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010001000: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8ce_ace_9bb_9bc_bdd_def_eff_eff_fff_eff_fff_fff_fff_eff_eff_dee_cee_abb_acd_9cd_8ce_7ce_7cf_7cf_7cf_7cf_8cf_8cf_7cf_8cf_8ce_def_eef_edf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dee_def_abc_acc_9cc_acd_acd_9cd_9bd_9cf_8cf_7cf_7df_6cf_6cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8be_ace_bce_cde_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_ffe_eee_cef_8ce_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_6cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010001001: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8df_7ce_9ce_dff_cee_eff_eff_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eff_fff_dff_cef_bff_8ce_8cf_8cf_8cf_7cf_8cf_8cf_8cf_8cf_9ce_def_eef_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_eff_eff_eff_eff_eff_eff_eff_dff_cef_9ce_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_9ce_def_cef_def_def_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_cff_8ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010001010: horiz=6144'h_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7be_9ce_9cd_dff_dee_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_eff_eff_dee_cef_acd_9cd_9be_9ce_8be_8cf_8cf_8ce_9ce_ace_eef_eef_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_eff_def_cdf_abd_ace_9ce_9df_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_9ce_def_def_def_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_cff_8cf_7cf_7cf_7cf_7cf_7ce_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7ce_7ce_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_7cf_7cf_7cf_7cf_7cf_8cf_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf;
				8'b010001011: horiz=6144'h_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_8ce_cef_cef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_eff_eff_cef_cef_8be_8ce_9df_9de_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_ffe_fff_fff_fff_fff_fff_fff_eff_dff_cff_cff_8ce_8cf_8cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_8ce_9cf_ace_eff_def_dee_eef_ddf_eef_eef_eef_eef_eef_eef_eef_eef_edf_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_fff_eff_def_cef_8ce_8cf_8cf_8cf_8cf_8ce_8df_7df_7cf_7cf_7cf_7cf_8cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7ce_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8df_7cf_7cf_7cf_7cf_7cf_8cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7ce_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf_7cf_8df_8df_7cf_7cf_7cf_7cf_7cf;
				8'b010001100: horiz=6144'h_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8cf_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8cf_8cf_8df_8cf_7cf_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_7cf_7cf_8cf_8cf_7cf_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_8df_8df_7cf_8ce_8bd_cef_def_eff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_def_def_9ce_9cf_8ce_9cd_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_cff_8bd_7ce_7cf_8cf_8cf_8cf_7cf_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7df_7cf_7ce_8cf_9ce_ace_bce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eff_eff_eff_fff_fff_fff_fff_fff_def_def_ace_9ce_9ce_9be_9cd_9cd_9ce_9df_7ce_7cf_7cf_7cf_8cf_7cf_8df_8df_7cf_7cf_7cf_7cf_8df_7cf_8cf_8cf_7cf_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8cf_8cf_8df_7df_7cf_7cf_7cf_7cf_8df_7cf_8df_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8df_7cf_7cf_7cf_7cf_8cf_8cf_7ce_8df_8df_7cf_7cf_7cf_7cf_8df_7cf_8cf_8cf_7cf_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7cf_7cf_8df;
				8'b010001101: horiz=6144'h_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_9df_8df_7ce_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_8ce_9de_9cd_def_def_dee_eee_eee_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_ffe_efe_fff_eff_dff_cef_9bd_9bd_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_fff_fff_fff_eff_eff_eff_eff_eff_eff_eff_eff_fff_eff_fff_eff_dff_9cd_8ce_8df_8df_8cf_7ce_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_8cf_9df_9ce_cff_def_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_eef_eff_def_def_dff_def_def_def_cef_cef_9ce_9cf_8cf_7ce_8df_8df_7ce_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_8cf_8df_8df_7ce_7ce_8df_8df_7ce_7ce_8df_8df_7ce_7ce_8df_8cf_8cf_8cf_8cf_8df_7ce_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df;
				8'b010001110: horiz=6144'h_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8cf_7cf_8cf_8cf_7cf_8cf_8cf_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8cf_7cf_8cf_8cf_7cf_8cf_8df_8cf_8cf_7cf_8df_7cf_8cf_8cf_8cf_8cf_8df_7ce_8cf_8cf_7cf_7cf_8df_8df_8cf_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8cf_8df_8ce_ade_ace_def_def_eef_ede_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_eff_eff_fff_fff_fff_def_cdf_bcd_abc_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eee_fff_fff_fff_eff_eff_eff_eff_fff_fff_fff_fff_eff_fff_fff_eff_eff_9cd_9ce_8df_8df_8df_7ce_8cf_8cf_7cf_8cf_8df_8df_8cf_7cf_8cf_8cf_7cf_7df_8df_8df_8df_7cf_7cf_7cf_8cf_8cf_8cf_9cd_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_def_dee_def_acd_9bc_9cd_8ce_8df_8df_7cf_7cf_8df_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8cf_7cf_8cf_8cf_7cf_7df_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8cf_7cf_7cf_7cf_8df_7cf_8ce_8ce_9df_9cd_9cd_8cd_9cd_9cd_9cd_9cd_9de_9cd_9cd_9cd_9ce_9df_8ce_8cf_8cf_8cf_8cf_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df_8df_8df_7cf_8cf_8cf_7cf_8cf_8df;
				8'b010001111: horiz=6144'h_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8cf_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8df_8df_7be_8cf_8cf_8df_8ce_8ce_8cf_8ce_8cf_7ce_8df_8cf_7ce_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7ce_8cf_8df_7cf_8cf_9df_9df_cff_cef_def_def_eef_eef_eef_eef_eee_eee_fff_fff_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_eee_eef_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_fff_fff_fff_eff_eff_eff_eff_fef_eee_eef_eef_eee_fff_fff_fff_ffe_ffe_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_cef_bef_8ce_7ce_8cf_8df_7cf_7ce_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_7cf_8df_7cf_7ce_8cf_8df_7cf_7cf_8df_8cf_8bd_9cd_def_def_edf_eef_eef_eef_eef_eef_eef_eef_eee_eee_fff_fff_fff_fff_fff_eff_def_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eee_eee_eee_eef_eef_eef_eef_eef_eef_eef_fff_dff_eff_fff_fff_eff_eff_cff_9ce_7ce_8df_8df_7ce_7ce_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7ce_8df_8df_7be_8ce_9ce_9ce_cff_dff_eff_eff_eff_eff_eff_eff_eff_fff_fff_eff_def_cef_8ce_9df_7ce_7cf_8df_8cf_7cf_7cf_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf;
				8'b010010000: horiz=6144'h_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_7cf_7cf_7cf_7cf_7cf_7cf_8cf_8cf_7ce_8cf_9cf_8cf_8df_8df_7cf_7cf_8cf_8df_8ce_9ce_9cd_acd_acd_acd_acd_acd_acd_9cd_9ce_8df_8df_7cf_8cf_8df_7ce_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_8cf_7cf_8cf_8df_8cf_7df_8df_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_eff_fff_fff_fff_fff_fff_efe_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eff_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dee_cef_8ce_7cf_7cf_7df_7df_7df_7df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8df_8df_7cf_7df_8df_8cd_acd_bcd_def_eef_eef_eef_def_eef_eef_dee_eee_eee_eef_eef_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eee_fff_fff_fff_fff_fff_fff_eff_def_acc_9de_8de_7ce_7cf_7cf_8df_8cf_8cf_7ce_7ce_8df_7cf_7cf_7df_7cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_7cf_7cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_7cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_8cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_7cf_8cf_8cf_9ce_9bc_acd_bdd_def_eff_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_dee_cdd_acc_add_9cd_9de_8ce_8cf_7cf_8cf_8df_8cf_8cf_8cf_8cf_7cf_8df_7cf_7df_7cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_7cf;
				8'b010010001: horiz=6144'h_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_8cf_8df_8df_7cf_7cf_8df_8cf_8ce_9ce_cff_cff_eff_eff_eff_dff_dff_eff_dff_cef_8bd_8ce_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_8cf_8df_7df_7ce_9ce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_fff_fff_eee_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_cff_8ce_8df_7ce_7ce_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7ce_8df_8cf_8cf_9ce_dff_def_def_eef_eef_eef_eef_eef_eef_eee_eee_eef_fff_fff_fff_fff_fff_ffe_ffe_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_eff_eff_fff_fff_fff_fff_efe_eff_eff_eff_cff_8cd_8cd_8cf_8df_8cf_7cf_8cf_8df_7cf_7cf_8df_8df_7cf_7ce_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7ce_8df_8df_8cf_7ce_8df_8df_7cf_7ce_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8cf_8df_8cf_7ce_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8cf_8ce_9ce_cff_def_eff_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_cff_bff_8bd_8ce_8df_8cf_7ce_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df_8df_8cf_7cf_8df;
				8'b010010010: horiz=6144'h_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8cf_7cf_8cf_8df_8df_7cf_8cf_7df_8df_7cf_8cf_8cf_8cf_8ce_9df_acd_acd_acd_def_eff_eff_fff_fff_eff_eff_eff_def_def_9bc_9cd_9ce_9df_8cf_7ce_7cf_8df_8cf_7cf_7df_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8cf_7cf_8cf_8df_8df_7cf_8cf_7df_8ce_9ce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_eff_eef_eee_eff_eff_fff_fff_eff_eff_fff_fff_eff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_8ce_8df_8df_7ce_7cf_8df_8df_7cf_8cf_8df_8cf_7cf_8cf_8df_8cf_7cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_9ce_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_ffe_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eee_eff_fff_eff_eff_fff_fff_fff_ffe_eff_eff_eff_dff_abd_acd_9cd_9ce_9cf_8cf_8cf_8cf_8cf_7cf_8cf_8df_8df_7ce_8cf_8df_8cf_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8cf_7ce_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8cf_7cf_8cf_8df_8df_7ce_8cf_8df_8df_7cf_8cf_8df_8cf_7cf_8cf_8df_8df_7cf_7cf_9ce_ace_abd_def_eee_eff_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_cef_9bc_9ce_9ce_9cf_8ce_8cf_8cf_8df_8cf_7cf_8cf_8df_8cf_7ce_8cf_8df_8cf_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf;
				8'b010010011: horiz=6144'h_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_8ce_8cf_8df_7cf_7ce_8cf_8df_7ce_7cf_8df_8cf_8ce_8ce_9df_9df_dff_def_eef_dee_eff_ffe_ffe_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_bff_9df_8ce_7ce_7ce_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_8df_8df_7cf_7ce_8df_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_dde_eee_fff_fff_eee_eee_fff_eff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dee_cef_8ce_7ce_8df_8df_7ce_7ce_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_9df_8cf_8cf_9cf_ace_dff_def_def_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_eff_eff_eff_eff_eff_eff_fff_fff_fff_fff_fff_eff_eef_fff_eff_def_def_cef_aef_8ce_8cf_8cf_8cf_7cf_7ce_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7ce_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_7df_8df_7cf_7cf_7cf_7cf_8df_7ce_8cf_8df_7cf_7ce_8cf_8df_7cf_7ce_8cf_8df_7cf_7cf_8cf_8df_7ce_abd_dff_def_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_dff_cef_cff_9ce_9cf_7cf_7cf_8cf_8cf_8df_7ce_8cf_8df_8cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_8cf_8df_7cf_7cf_8cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf_7cf_7cf_8df_7cf;
				8'b010010100: horiz=6144'h_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_8cf_8df_7cf_7cf_7cf_8cf_8df_8df_7cf_7cf_8df_8ce_7bd_8ce_9ce_9bd_ace_ace_bde_def_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_cff_9ce_8ce_7ce_7cf_8df_7cf_7df_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_7cf_7cf_8df_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eef_fff_eff_eef_eef_eff_eff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_eff_eff_fff_fff_fff_fff_eff_fff_eff_eef_def_cef_8ce_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_8cf_8df_8cf_8cf_7cf_7cf_8df_8df_8cf_8cf_9df_cef_cef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eff_efe_fff_fff_fff_fff_fff_eef_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eee_eef_def_cdf_ace_8ce_9ce_8cf_7ce_7ce_7cf_7cf_8df_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_7cf_8df_7cf_8cf_8cf_8df_7cf_7cf_7df_8df_7cf_8cf_7cf_8df_7cf_6cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_7cf_8cf_8cf_8cf_9df_bcd_eff_def_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_def_acd_adf_8ce_7cf_8cf_8df_7cf_7cf_7cf_8cf_8df_7cf_8df_8cf_7cf_8cf_8df_8cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_8cf_8df_8cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf_7cf_7cf_8df_8df_7cf_8df_7cf_8cf;
				8'b010010101: horiz=6144'h_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7ce_8ce_9cf_9cc_cef_cef_def_eff_def_eef_ede_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_dff_8bd_8ce_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7ce_7ce_8df_7df_7ce_9ce_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_fff_fff_eef_eef_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_eef_dee_eef_eff_eff_fff_fff_fff_eff_def_eef_def_cef_9df_8df_7cf_7ce_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7ce_8df_7cf_7cf_8ce_9ce_abd_eff_def_fef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eee_eef_eef_eef_eef_cef_cef_bef_8cd_9df_8cf_7cf_7cf_8df_8cf_7cf_8df_8df_7cf_8cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7ce_8df_8df_7cf_7cf_8df_9df_8ce_8ce_8df_8df_8ce_8ce_9df_9df_8ce_7cf_7cf_8cf_7ce_7ce_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_8ce_9ce_dff_eef_def_eef_def_def_def_def_def_eef_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_eff_eff_eff_eff_eff_fff_fff_fff_fff_eff_dff_cef_9ce_8cf_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8cf_8df_7cf_8cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_8cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df_8df_7cf_7cf_8df;
				8'b010010110: horiz=6144'h_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8df_8df_7cf_8cf_8ce_9df_8bd_ace_bcd_def_eef_eef_eef_eef_eee_eee_eef_eef_dee_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_eff_9bc_9ce_8cf_8cf_8cf_8cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8df_8cf_7ce_8df_7df_8cf_9be_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_eee_eef_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eff_fff_fff_fff_eff_def_eff_def_bef_9df_8df_8df_7ce_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_7cf_7cf_8cf_8ce_acd_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_fff_eff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eef_eef_eef_eef_eef_eef_dee_def_acd_9ce_9ce_8ce_7be_8df_8df_7cf_8cf_8cf_8cf_8cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8cf_7cf_8cf_8cf_8cf_7cf_8df_8cf_8cf_8ce_9de_9cd_9cd_9cd_9cd_9cd_9cd_9cd_acd_9cd_9cd_8ce_7ce_8cf_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_7cf_8cf_8cf_9ce_acd_def_eef_eef_eef_def_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_cef_ade_9df_8ce_8ce_8df_8df_8df_7cf_8cf_8df_8cf_7cf_7cf_8cf_8cf_8cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_8cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df_8df_8df_7cf_8cf_8cf_8cf_7cf_8df;
				8'b010010111: horiz=6144'h_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_8cf_8df_7cf_7cf_7ce_8cf_8df_8ce_9ce_cef_cef_def_def_dde_eef_eef_eef_eef_eef_eef_eee_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_eff_dff_bef_8cf_8cf_8df_8cf_8cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_8cf_8df_8cf_7cf_7cf_8df_9ce_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_dee_def_def_def_ace_9ce_8df_7ce_8df_8df_7ce_8cf_8df_8cf_7cf_7cf_8cf_8df_7cf_8cf_8df_8cf_8cf_7cf_8cf_9df_7ce_7cf_8df_8cf_8ce_9cd_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eee_eee_eee_eee_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eee_eee_eee_eee_eef_eef_eee_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_def_def_eef_eef_eee_fde_fdf_fef_eef_cef_cef_bef_8cd_7cf_7cf_8df_7cf_8cf_8df_8cf_8cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_8df_7ce_8ce_9df_ace_dff_dff_eff_eff_eff_eff_eff_eff_eff_eff_cef_bef_8bd_8cf_8df_8cf_8cf_8cf_8df_8cf_8cf_8bf_8cf_8df_8cf_9ce_cff_eff_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_ffe_fff_fff_eff_dff_cff_9ce_8ce_8ce_7ce_8df_8cf_8ce_7cf_8df_8cf_7cf_8cf_8df_8cf_8cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_8cf_8df_8cf_8cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf_7cf_8cf_8df_7cf_7cf_8df_7cf_7cf;
				8'b010011000: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8df_8cf_8cf_8cf_8df_8df_7cf_7df_8df_9ce_ace_acd_cde_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_eff_fff_fff_fff_eee_cef_9ce_8cf_8cf_8cf_8cf_7cf_8df_8cf_8cf_8cf_8cf_8cf_7cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_7cf_8cf_8cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_7cf_8cf_8cf_7cf_8cf_8df_8cf_8cf_7cf_8cf_8cf_7cf_7cf_7df_9df_bef_cdf_def_eef_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eee_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_eee_eee_eee_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_bcd_ade_8ce_7cf_8df_7cf_7cf_7cf_8cf_8cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_9ce_cef_cdf_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_def_dff_cef_bef_8ce_8cf_8df_8cf_8cf_7cf_8cf_8cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_7cf_8cf_9ce_9cd_abc_acc_bcc_dee_eff_eff_fff_fff_efe_eff_eff_eff_eff_dee_dee_abc_acd_acd_9de_7ce_8df_7df_8df_7ce_8cf_8df_8cf_8ce_9cd_def_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_eff_eee_cee_acc_acd_acc_acd_ace_ade_9cd_8de_8df_7cf_7ce_7cf_7cf_8df_7ce_8cf_8df_8cf_8cf_7cf_8cf_8cf_7cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8df_7cf_7cf_7cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7cf_8cf_8df_7ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010011001: horiz=6144'h_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7cf_8cf_8df_8cf_8df_8df_8df_7df_8cf_9ce_cef_cdf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_fff_fff_fff_fff_fff_eff_eff_eff_fff_fff_fff_eff_dff_9ce_8df_8df_8df_8df_8df_7cf_7cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8df_8df_8df_8df_7df_7cf_8ce_9ce_9cd_def_def_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cff_9df_8df_7cf_7cf_8cf_8df_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_9ce_8bd_9bd_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_dee_def_eef_eef_eef_eef_def_eef_eef_eef_def_cef_9cd_9cf_9df_8df_7ce_8cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7cf_7cf_8df_8df_8ce_ade_dff_def_eff_eff_eff_eff_fff_eff_fff_fff_fff_eff_eff_eff_fff_eff_fff_eff_def_cef_9ce_9df_9df_8cf_8cf_8df_8cf_8ce_9de_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_eff_fff_eff_eff_eff_eff_dff_cef_bff_8cd_8ce_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8df_8df_8df_8df_8df_7cf_8cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8df_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df_8df_7ce_8cf_8df_8cf_8df_8df_8df;
				8'b010011010: horiz=6144'h_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_8ce_9be_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_fff_fff_eff_eff_fff_fff_fff_eff_eff_dff_8ce_8df_8df_8df_8df_8de_8de_7ce_7df_8df_8df_8cf_9df_8cf_8cf_7cf_8df_8df_8df_8cf_8df_8cf_8cf_7cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_7cf_8df_8df_8df_8df_8df_8cf_8cf_7cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8ce_ade_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cef_9ce_8df_8df_7cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_7ce_8ce_bef_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_eef_dee_def_eef_eef_eef_def_eff_def_def_cef_bef_9ce_8cf_9df_8cf_8cf_7cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_7cf_7cf_8df_8ce_9de_acd_dff_eee_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_def_acd_ace_ace_9cf_9cf_8cf_8cf_8ce_ade_bce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_dfe_cef_9bd_9cd_9ce_adf_8cf_8cf_8df_8cf_8cf_7cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8df_8cf_8df_8cf_8cf_7cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df;
				8'b010011011: horiz=6144'h_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8cf_8cf_8df_8cf_8df_8df_8df_9df_9ce_ace_def_def_dee_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_edf_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_eff_fff_fff_fff_eff_dee_cef_9ce_9ce_8cf_8cf_9ce_9de_9df_8ce_8df_8df_8df_8df_8cf_8df_8df_8df_8df_8df_8df_8cf_8cf_8df_8df_8cf_8df_8df_8df_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8df_8cf_8cf_8df_8df_8cf_8df_8df_8df_8cf_8cf_9df_8cf_8df_8cf_9ce_9ce_bce_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_cef_9ce_8df_8df_8df_8cf_8df_8df_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8df_8cf_8df_8df_8df_8ce_8ce_9ce_cef_def_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_eef_def_def_cff_9ce_9ce_9ce_9ce_9df_8df_8df_8df_8df_8cf_8df_8df_8df_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9df_cef_cef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_cef_ace_8df_9df_ace_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_eff_fff_eff_cef_cef_9ce_8cf_8df_8df_8df_8cf_8df_8df_8df_8cf_8cf_8df_8df_8cf_8df_8df_8df_8cf_8cf_8df_8df_8cf_8df_8cf_8df_8cf_8df_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf;
				8'b010011100: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9ce_ace_bde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_eff_eff_fff_fff_fff_fff_eef_eef_def_ace_ace_ace_ace_ace_ace_ace_9cf_8cf_8df_7df_8df_8cf_8df_8df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8ce_9ce_bce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_dee_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_cdf_ace_9df_8cf_8df_8cf_7cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8cf_8cf_8cf_8df_8ce_bef_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_def_eef_eef_def_cef_aef_9ce_9cf_8cf_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_7df_8df_8df_9ce_9ce_cef_def_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_ffe_fff_eef_cef_ace_9df_8cd_acd_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_eff_def_dff_9ce_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010011101: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_9ce_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_ede_eef_eef_def_def_def_def_def_def_cef_9ce_9df_8df_8df_7df_8df_8df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9cf_cef_cdf_ddf_dde_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_dff_bef_9ce_8ce_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_9cf_9cf_8cf_8cf_9df_9ce_ace_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_def_ddf_ddf_ddf_cdf_acd_9ce_8ce_9df_8cf_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_9ce_acd_def_def_eef_eee_eee_eee_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_ffe_ffe_ffe_fff_eff_dff_bef_acd_acd_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eee_eee_fff_fff_fff_fff_fff_fff_eff_eff_eff_eff_eff_fff_efe_fff_eff_dff_9cd_9df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010011110: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_8cf_8ce_acd_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_def_eef_dee_def_def_abc_acd_ade_9de_8ce_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9cf_cef_cdf_ddf_dde_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_def_cef_abd_ace_9ce_9df_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_9df_ace_ace_def_def_def_def_def_def_def_def_def_ddf_eef_def_eef_eef_eef_eef_eef_def_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_ddf_ddf_ddf_cdf_ade_9de_8ce_8cf_8df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_9ce_ade_bce_def_eef_eef_eee_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_fff_fff_eef_def_bce_bcd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eee_eee_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_eff_eff_efe_fff_eff_eff_acd_9de_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8df_8df_8df_8ce_8ce_9de_9ce_9ce_9ce_9ce_9df_9df_8ce_9df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010011111: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8cf_8cf_9ce_9cd_def_eef_ede_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_eff_def_eef_eef_eef_eef_eef_eef_ddf_def_dee_eee_eee_eee_eee_eef_eef_eef_eef_eef_eef_fff_eff_eff_efe_fff_eff_eff_dff_9ce_8df_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_9cf_9cf_cef_cdf_dde_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_def_def_eef_eef_eef_def_eee_eee_def_cef_bef_9ce_9cf_9ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_9cf_8be_def_def_ddf_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_ddf_def_dde_def_def_def_def_def_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_ddf_ddf_ddf_def_cff_bef_8ce_9cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_adf_cef_cef_def_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_eff_fff_fff_eff_eff_fff_fff_fff_fff_eff_fff_fff_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_fff_fff_fff_eff_eff_eff_eff_eef_eee_eef_eee_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_ffe_eff_def_bef_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8df_8df_8ce_8ce_9ce_dff_def_def_def_cef_bef_8ce_8ce_9df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100000: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8ce_bde_bcd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_ffe_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eff_fff_fff_fff_ffe_ffe_ffe_eff_dfe_bcd_bdf_9ce_8ce_8cf_7df_8df_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9df_bef_bdf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_dee_eff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_dee_eff_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_cde_abd_ace_ace_adf_9cf_8ce_8df_8df_8df_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_9cf_9ce_cef_ddf_edf_ddf_def_ddf_ddf_ddf_ddf_ddf_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_def_def_ddf_ddf_def_def_def_dee_cef_acd_ace_9ce_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_9ce_def_def_def_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_eff_fff_fff_fff_fff_fff_efe_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eff_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_efe_efe_dfe_cff_9ce_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8df_8df_8df_8df_8df_9ce_ade_bce_eef_fef_eef_eef_def_bef_9cd_acd_9cc_9cd_9ce_9df_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100001: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_adf_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_ffe_ffe_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_ffe_ffe_efe_eff_eff_dff_9ce_9ce_8ce_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9df_9cd_acd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_fff_fff_fff_fff_eff_fff_fff_fff_fff_eff_fff_eff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_cef_bef_9ce_8ce_8df_8df_9cf_9df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_9cf_9ce_cef_def_edf_def_def_def_def_def_def_def_def_ddf_ddf_def_def_def_def_def_ddf_def_def_def_def_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_cef_cef_cef_cef_cef_adf_8ce_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_9ce_def_def_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_fff_fff_eee_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_9ce_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8ce_9ce_ace_dff_def_eef_eef_eef_eef_eef_def_eef_def_eef_def_cef_bef_9ce_8df_8df_8cf_8cf_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100010: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9cf_ace_dff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_ffe_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_eff_fff_fff_fff_fff_efe_eff_eff_dff_acd_acd_ace_ade_9cf_9df_8ce_8df_8df_8cf_8cf_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8cf_9ce_ace_bce_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_bdf_ace_9ce_ade_adf_9ce_9df_8ce_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9cf_bef_cdf_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_cef_cef_cef_cef_cef_cef_bef_bef_adf_8cf_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9cf_ace_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_eff_eef_eee_eff_eff_fff_fff_eff_eff_fff_fff_eff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_9cf_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8ce_9ce_9ce_ace_bce_def_eef_def_eef_eef_eef_eef_fdf_fdf_fef_fef_eef_ddf_cef_bce_9df_8df_8cf_8df_8df_8df_8df_7df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100011: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9df_ace_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_ffe_eff_eff_fff_fff_fff_fff_fff_eff_eff_eff_eff_def_dff_cef_bef_9cd_9cf_9df_8cf_8cf_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_9ce_ade_dff_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eef_eee_eee_eee_eee_eef_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_def_cef_cdf_def_def_cef_bef_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8cf_9cf_9be_ace_def_cef_def_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_ddf_cdf_bef_9ce_9ce_9ce_9cf_9cf_9ce_8ce_8cf_9df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9cf_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_dde_eee_fff_fff_eee_eee_fff_eff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_fff_eff_eff_eff_eff_eff_fff_fff_fff_fff_def_cef_9ce_8df_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_9ce_cef_cef_def_eef_def_def_def_eef_eef_eef_eef_fef_eef_eef_eef_dee_def_dff_dff_cff_9ce_9ce_9cf_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100100: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_8df_adf_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eff_eff_fff_fff_fff_fff_fff_eef_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eef_eef_def_cde_acd_9df_9cf_9cf_9cf_8ce_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8ce_9ce_bce_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_def_def_def_def_cdf_bdf_ade_9df_8ce_8df_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_9cf_9cf_bef_cef_cdf_cdf_def_def_ddf_ddf_def_def_cdf_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bdf_bdf_cdf_cef_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_cdf_cef_cef_adf_8ce_8df_8df_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9cf_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eef_fff_eff_eef_eef_eff_eff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_eff_eff_eff_eff_eff_eff_eff_fff_fff_fef_eef_cef_9df_8ce_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_9cf_9ce_cef_cef_def_eef_eef_def_eef_def_def_eef_eef_def_def_def_def_dee_def_def_def_cef_ace_ace_ace_9cf_9cf_9df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100101: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8ce_9ce_acd_def_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_eff_efe_fff_eef_eef_eef_eef_def_dff_dff_cef_9bd_9ce_9cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9cf_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eee_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_ddf_def_def_cef_def_9bc_acd_bff_bef_8ce_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8ce_9cf_9bd_9cd_abd_def_def_def_def_def_bef_9ce_9ce_9ce_9de_9df_9df_9df_9ce_9ce_9ce_9ce_8ce_9ce_9ce_bef_def_def_def_def_def_def_def_def_def_def_def_def_def_cef_cef_9bd_9ce_9ce_8ce_8df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_9cf_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_fff_fff_eef_eef_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_def_eef_dee_def_def_def_def_dee_dee_def_def_eef_def_cef_9ce_9ce_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_9cf_9ce_bef_cef_def_ddf_dde_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_def_def_def_ddf_cdf_def_cef_cef_cef_9ce_9ce_9df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100110: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8cf_9cf_9cd_dff_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_fff_eff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eef_eef_eef_eef_eef_def_def_def_acd_ace_9ce_9ce_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_9ce_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_eef_eff_eff_fff_fff_fff_fff_eff_fff_eff_fff_eef_def_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_def_def_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_ddf_def_def_cef_cdf_bce_ace_bef_aef_9ce_8ce_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_9df_8ce_9df_bef_cef_cef_cef_cef_adf_9ce_9ce_9df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8ce_9df_aef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bef_bef_adf_9cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_ace_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_eee_eef_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_ade_ace_9ce_9ce_8ce_8cf_8df_8df_8df_8df_8df_8cf_8cf_9df_bef_cef_cef_cdf_def_def_ddf_def_def_def_def_edf_ddf_ddf_def_def_def_cef_def_cef_bef_cef_bef_aef_9ce_8ce_9df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010100111: horiz=6144'h_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_9cf_9cd_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eef_eee_eee_eee_eee_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eee_eee_eef_eef_eef_eef_eee_eee_eef_fff_fff_fff_fff_fff_eff_eff_eff_def_def_eef_eef_fef_eee_eef_eef_def_cef_cef_bef_8cd_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_ace_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_dee_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_ddf_def_def_def_eef_def_eef_eef_eef_eef_eef_eef_ddf_ddf_def_ddf_cdf_bdf_9cd_ace_cff_cef_9ce_9ce_9ce_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_7df_8ce_8ce_9de_9ce_9ce_9ce_9cf_9cf_8cf_9df_8df_8df_8df_8df_8df_8df_8df_8df_8df_8cf_8cf_8ce_9cf_9cf_9cf_9cf_9cf_9cf_9cf_9cf_9ce_9ce_9ce_9ce_8ce_8ce_8ce_8df_8df_8df_8df_8cf_8cf_8cf_8df_8df_8df_8df_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8df_8cf_9ce_cef_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eef_eef_def_cef_bef_8ce_8cf_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8ce_9ce_9ce_acd_cef_def_ddf_ddf_ddf_def_cef_ddf_ddf_def_cef_cef_9ce_8ce_9df_9cf_9cf_9cf_8ce_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf;
				8'b010101000: horiz=6144'h_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8df_8df_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8df_8df_9df_bff_bdf_eef_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_eff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_bdf_bef_9df_8df_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8cf_8cf_9ce_def_eef_eef_eef_def_def_def_def_def_def_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_ddf_def_ddf_def_def_def_eef_eef_eef_eef_eef_eef_def_def_cef_bef_bef_bdf_9ce_9df_aef_aef_9de_7df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8cf_8ce_ade_acd_add_acd_acd_acd_acd_ace_9ce_9cf_8cf_8df_8df_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8cf_8df_8df_8cf_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8cf_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8df_8df_8df_8cf_9cf_cef_cdf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eee_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_eee_eee_eee_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fef_eef_def_cef_bef_cff_aef_8ce_8cf_8cf_8df_8df_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_ace_bef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_aef_9cf_9cf_9cf_8cf_8df_8df_8cf_8df_8df_8df_8df_8cf_8df_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf;
				8'b010101001: horiz=6144'h_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_9df_9ce_9cd_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_acd_9ce_9df_8df_8df_8cf_8df_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8df_8df_8df_8df_8cf_ace_def_eef_eef_eef_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_def_ddf_ddf_ddf_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_cef_9bd_9ce_9ce_9ce_9cf_8ce_8ce_8ce_8df_8df_8df_8df_8cf_8cf_8cf_8cf_8df_8cf_8cf_8df_8cf_8df_8df_8df_8cf_8df_8cf_8cf_9ce_9ce_cef_def_dff_eff_eff_eff_eff_eff_cef_cef_ace_8de_8df_8cf_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8df_8df_8df_8df_8df_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_8df_8df_8cf_9ce_acd_def_def_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_cef_9bd_9ce_8ce_9ce_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8cf_8cf_8cf_8cf_8cf_9ce_9ce_9ce_8bd_9ce_9ce_9ce_9ce_9ce_9ce_9ce_9ce_8ce_9cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_8df_8df_8cf_8cf_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf;
				8'b010101010: horiz=6144'h_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_9df_9cf_9ce_cef_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_bde_9ce_8ce_8df_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_9cf_ace_def_eef_eef_eef_ddf_def_def_def_def_def_def_def_def_def_def_def_def_ddf_eef_eef_eef_def_def_def_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_eef_def_eef_eef_eef_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_ddf_def_def_ddf_ddf_ddf_def_def_def_def_def_def_eef_eef_eef_eef_def_def_acd_ade_9ce_9ce_9cf_9df_8cf_8cf_9df_8cf_8df_9df_8cf_8cf_8cf_8cf_8cf_7df_8df_8df_8cf_8df_8df_8cf_8df_9be_ace_ace_ace_acd_def_def_eee_fff_fff_fff_fff_fff_def_def_acd_ace_9ce_9ce_8ce_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8df_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8df_8df_8cf_8df_8df_8df_8df_8df_8df_8df_8ce_9ce_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cef_9cd_8ce_9df_8cf_8cf_8cf_8df_8cf_8cf_8cf_8df_8df_8cf_8cf_8cf_8cf_8cf_8cf_9df_8cf_8cf_8cf_8cf_8cf_8cf_8ce_8ce_8df_8cf_8df_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8df_8df_8df_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf_8cf_8cf_8df_8cf_8cf_8cf_8cf_8cf;
				8'b010101011: horiz=6144'h_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8df_8df_8df_9df_9df_8cf_8df_8df_8df_8df_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8ce_9df_9df_8bd_9cd_def_def_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_eef_def_def_eef_fff_fff_fff_eff_dff_cff_9de_8cf_9df_9df_8cf_8cf_8cf_8df_8df_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8df_8ce_adf_bde_def_eef_edf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_def_ddf_ddf_def_def_def_def_ddf_def_ddf_eef_eef_eef_eef_def_def_cef_cef_bdf_ade_bef_bef_9ce_8cf_9df_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8df_8df_9df_8ce_8ce_9ce_9ce_9ce_abd_def_def_def_eef_fff_fff_ffe_fff_fff_fff_fff_ffe_ffe_fff_eff_eff_cef_bef_8ce_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8df_8df_8df_8df_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8df_9de_9ce_ace_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cef_9ce_9df_aef_9df_8df_8df_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8df_9ef_8df_8cf_8cf_8cf_8cf_8cf_8df_9df_8df_8cf_8df_8df_8df_8df_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf_8cf_9df_9df_8cf_8cf_8cf_8cf_8cf;
				8'b010101100: horiz=6144'h_8df_9df_9df_8ce_8df_8cf_8cf_8cf_9df_9df_9df_8ce_9df_8cf_8cf_8cf_9df_9df_9df_8cf_8cf_8cf_8cf_8cf_9df_9df_9df_8cf_8cf_8cf_8cf_8cf_9df_9df_9df_8cf_8df_8df_8cf_8cf_8df_9df_9df_8ce_8cf_8cf_8df_8df_9df_9df_9df_9df_8df_8cf_8df_8cf_9df_9df_9df_8cf_9df_8cf_8cf_8cf_8df_9df_9df_8ce_8df_8cf_8cf_8cf_8df_9df_9df_8cf_8df_8cf_8cf_8cf_9cf_9df_9df_8ce_9de_bef_def_eef_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_eef_def_eff_eff_fff_fff_fff_eff_def_cff_9ce_9cf_9df_9df_8cf_9df_8cf_8cf_8cf_8df_9df_9df_8cf_8df_8df_8cf_8cf_9df_9df_9df_8cf_8cf_8cf_8cf_8cf_9df_9df_9df_8cf_8df_8cf_8cf_8cf_9df_9de_ade_cef_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_def_def_def_def_def_ddf_ddf_def_def_def_eef_def_eef_eef_eef_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_ddf_def_def_def_eef_eef_eef_eef_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_eef_eef_eef_def_def_def_cef_bcd_bde_cef_cef_ace_ade_9ce_9df_9df_8df_8df_8df_8df_8cf_8cf_9df_9df_9cf_adf_ace_ace_ace_ace_bce_def_def_eef_eef_fff_fff_ffe_fff_fff_fff_fff_fff_fff_fff_fff_eff_def_cff_9ce_8ce_8df_8cf_8cf_8ce_9df_9df_8ce_8cf_8df_8cf_8cf_9cf_9df_9df_8cf_8df_8df_8df_8cf_8cf_9df_9df_8cf_8df_8cf_8cf_8cf_8df_9df_9df_8ce_8df_8cf_8cf_8cf_9df_9df_8df_8df_8df_8cf_8cf_8cf_8df_9df_9df_8ce_8df_8cf_8cf_8cf_9cf_9df_9df_8ce_8ce_ace_bdf_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_dee_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_cdf_ace_9df_9df_9df_8cf_8cf_8cf_8cf_8cf_9df_9df_8df_8cf_8df_8cf_8cf_8cf_8cf_9df_9df_8ce_8df_8cf_8cf_8cf_8df_9df_9df_8cf_8df_8cf_8cf_8cf_9cf_9df_9df_8cf_9df_8cf_8cf_8cf_8df_9df_9df_8cf_8df_8cf_8cf_8cf_8df_9df_9df_8ce_8df_8cf_8cf_8cf;
				8'b010101101: horiz=6144'h_9df_8ce_8df_9df_9df_8df_9df_9df_9df_8ce_8df_9df_9df_8df_9df_9df_9df_8ce_8cf_aef_9df_8df_9df_9df_9df_8ce_8cf_9df_9df_8df_9df_9df_9df_8ce_8cf_aef_9df_9df_9df_9df_9df_8ce_8cf_9df_9df_8cf_8df_9df_9df_8ce_9df_9df_9df_8df_9df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8ce_8df_9df_9df_8df_9df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8ce_8df_9ef_9df_9ce_bce_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_def_def_eff_fff_fff_fff_fff_fff_eff_dff_ade_9df_9ce_9cf_9df_9df_8cf_9df_9df_9df_8ce_8cf_9df_9df_8df_9df_9df_9df_8ce_8cf_aef_9df_8df_9df_9df_9df_8ce_8cf_9df_9df_8df_9df_9df_9df_8ce_9ce_cef_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_dde_def_def_def_ddf_def_def_def_def_def_def_cef_def_bef_9ce_8df_9df_9ef_8df_9df_9df_adf_ace_ace_def_def_def_def_def_eef_def_eef_eef_eee_fff_fff_ffe_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_ade_9df_9df_8df_9df_9df_8ce_9df_9df_9df_8df_8df_9df_9df_8ce_9df_9df_9df_8df_9df_8df_9df_8cf_8cf_9df_9df_8df_9df_9df_9df_8ce_8df_9df_9df_8cf_9df_9df_9df_8ce_8cf_aef_9df_8cf_9df_9df_9df_8ce_8df_9df_9df_8df_9df_9df_adf_8ce_9df_9df_adf_cef_def_ddf_dee_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_dff_cff_9ce_9ce_adf_9df_9cf_9df_9df_9df_8cf_8cf_9df_9df_8df_9df_9df_9df_8ce_9df_9df_9df_9cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9cf_9df_9df_8cf_9df_9df_9df_8ce_8df_9df_9df_8df_9df_9df_9df_8ce_8df_9df_9df_8df_9df_9df;
				8'b010101110: horiz=6144'h_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_8df_8cf_9df_9df_8cf_9df_9df_9df_9cf_9cf_9df_9df_8ce_9df_9df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_9cf_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8ce_9df_9df_adf_ace_def_def_def_def_def_def_def_def_def_ddf_eef_def_eef_eef_eef_eef_eef_def_def_eef_eef_eef_eef_eef_ddf_def_def_def_def_ddf_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_ddf_def_ddf_def_eff_eff_fff_fff_ffe_fff_eff_eff_bde_adf_9ce_9ce_9df_9df_9df_9df_9df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_8df_9ce_bef_cdf_def_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_ddf_def_ddf_def_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_cef_ace_9ce_9df_8df_9df_9ce_adf_bde_bce_bde_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_fff_eff_eff_bde_bdf_9ce_9df_9ce_9df_8cf_8ce_9df_9df_8cf_9df_9df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_8cf_8ce_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_9cf_8ce_adf_adf_cef_def_ddf_dee_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cef_acd_acd_adf_adf_9cf_9cf_9df_9df_9cf_8cf_9df_9df_9df_9df_8df_9df_9df_8ce_9df_9df_9df_9df_9df_9df_9cf_8ce_9df_9df_9df_9df_9df_9df_9cf_8ce_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_8df_9df_9df_8cf_9df_9df_9df_9df_8df;
				8'b010101111: horiz=6144'h_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_9ce_9cf_adf_9df_8ce_9cf_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_9ce_cef_cef_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_dde_dde_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_ddf_def_ddf_def_dee_dde_fff_fff_ffe_fff_fff_eff_dff_cff_ade_9de_9de_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8df_9df_9df_9bd_9cd_cef_def_cdf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_cef_cef_def_def_def_def_ddf_ddf_def_cdf_def_def_def_ddf_ddf_ddf_ddf_def_cef_8bd_9df_adf_adf_cef_def_dff_def_eef_eef_eef_eef_eef_edf_edf_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_fff_dee_eff_eef_def_def_bef_9cd_8ce_adf_9df_8ce_8cf_9df_9df_8cf_8ce_9df_9df_8cf_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9ef_9df_8ce_ace_cef_cef_dee_dee_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_def_def_cef_cef_adf_9df_9df_8cf_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8cf_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce;
				8'b010110000: horiz=6144'h_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_8df_8df_9df_9df_9df_9df_8df_8df_8df_8df_9df_9df_9df_8df_8cf_9df_9df_8ce_9df_9df_8cf_9cf_9df_9df_9cf_ade_acd_bde_bdd_acd_acd_bde_bde_ace_ade_9df_9df_8cf_9cf_9df_9df_8cf_9df_9df_9df_8df_9df_9df_9df_9cf_9df_9df_9df_9cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8df_9df_9df_9df_8df_9df_9df_9df_9ce_ace_cef_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_def_def_ddf_def_def_ddf_ddf_def_fff_eff_eff_fff_eff_eff_eef_dff_ace_9df_9df_9df_9df_9ce_9df_8df_9df_9df_8cf_8cf_9df_9df_8cf_9df_9df_9df_8ce_9df_9df_8df_8df_9df_9df_9df_8ce_9df_9df_9df_8ce_8df_8df_8df_8cf_9df_bef_bef_bef_cde_def_def_ddf_ddf_ddf_eef_ddf_def_def_def_dde_ddf_def_def_def_cef_def_def_def_ddf_def_ddf_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_cdf_bef_bef_cdf_cef_def_dde_eef_dde_def_cef_def_def_def_def_def_def_def_def_def_def_def_def_dee_def_def_def_ddf_def_eef_dde_dde_def_def_cef_cef_bef_bdf_cef_cef_bef_bdf_cef_cef_bef_bdf_cef_cef_bef_bdf_cef_bef_bef_aef_9ce_ade_ade_bde_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fef_eef_eef_eef_eef_def_cde_bcd_ace_bce_bce_9ce_9df_9df_9df_7cf_8cf_9df_9df_8ce_9df_9df_8df_8df_9df_9df_9df_8cf_8df_8ef_8cf_8df_8df_9df_8df_7ce_8df_9df_9df_8cf_8df_9df_8df_8cf_9df_9df_9df_9ce_9df_9df_9df_8df_9df_9df_9df_8df_9df_9df_9df_9df_9cf_bef_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_dee_eff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_dee_eff_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_bce_bde_ace_adf_adf_9de_8df_8df_9df_9df_9cf_8df_9df_9df_8cf_9df_9df_9df_8df_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf;
				8'b010110001: horiz=6144'h_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_9df_9df_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8cf_9cf_adf_9df_8ce_8df_adf_9df_9cf_ace_cff_def_eff_eff_eff_eff_eff_eff_dff_cff_9cd_9ce_aef_9df_8ce_9df_9df_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_ace_cef_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_def_def_ddf_def_dee_fff_fff_eff_fff_eff_cff_9cd_8cf_9df_9df_8ce_8cf_9df_9df_8ce_8df_9df_9df_8ce_8cf_9df_9df_8ce_8cf_9df_9df_8ce_8cf_9ef_9df_8ce_8df_9df_9df_8ce_8df_9df_9df_8cf_8cf_aef_9df_8ce_9ce_ade_bde_cef_def_def_ddf_ddf_def_ddf_ddf_ddf_def_ddf_ddf_ddf_def_def_def_def_def_ddf_def_def_ddf_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_def_def_cdf_9bd_9ce_adf_ade_cef_def_def_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_def_ddf_def_ddf_def_ddf_def_def_cef_ace_9cf_9ce_9ce_adf_9cf_9ce_9ce_adf_adf_9ce_9ce_9df_adf_9ce_9ce_adf_9cf_9ce_9ce_adf_ade_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_fff_fff_fff_fff_fff_fff_fff_eff_dee_eef_eef_eee_eef_def_eef_eef_eef_def_def_def_cef_cef_9ce_8ce_9df_9df_8cf_9cf_adf_9df_8ce_8cf_9ef_9df_8ce_9df_9df_9df_8cf_8df_adf_9df_8ce_8ce_9df_9ef_8ce_8ce_9df_9df_8cf_8cf_9ef_9df_8ce_9cf_adf_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_9df_adf_ace_bce_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_fff_fff_fff_fff_eff_fff_fff_fff_fff_eff_fff_eff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_dff_cef_bef_9ce_9ce_9df_aef_8ce_9df_9df_9df_8cf_8cf_9df_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef_9df_8ce_8cf_aef;
				8'b010110010: horiz=6144'h_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_9df_9cf_9df_9df_9df_8cf_9df_8df_8df_8cf_9df_9df_8ce_9de_adf_bce_acd_bcd_def_eef_eff_fff_fff_eff_eff_fff_eff_cee_acd_acd_bde_adf_8ce_9df_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_adf_cef_cdf_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_dee_eef_fff_fff_eff_eff_eff_cff_9ce_9cf_8df_8df_8cf_8df_9df_9df_9de_8ce_9df_9df_9df_9cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9cf_9df_9cf_bdf_cef_cef_cef_cef_cef_cef_cef_cdf_def_def_ddf_ddf_ddf_ddf_ddf_def_cdf_cef_cdf_cdf_def_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_cdf_cde_cef_cef_cef_bdf_ace_9ce_adf_aef_bff_cff_cef_cdf_cdf_cdf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_cdf_cef_cef_cef_cef_cef_cef_bef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9de_9df_9df_9cf_9df_9ce_adf_ade_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eff_fff_fff_fff_fff_fff_fff_eff_eef_eef_eee_eef_eef_eef_eef_def_eef_def_eef_eef_ddf_def_ace_9ce_9df_9df_8df_8ce_aef_9df_9df_9cf_9df_8df_8df_9df_9df_9df_8cf_9ce_adf_ade_ace_acd_bde_ade_9ce_9ce_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_8df_8df_9df_adf_bdf_bcd_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_cef_bdf_acd_acd_ace_ade_9ce_adf_9df_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df;
				8'b010110011: horiz=6144'h_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_9df_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8df_9df_9df_9ce_9ce_adf_adf_dff_eef_eef_dee_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_def_bff_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_9ce_ace_ace_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_ddf_def_ddf_def_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_def_cff_adf_9cf_8cf_9df_adf_9df_8ce_9df_9df_9df_8ce_9df_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_9ce_adf_adf_9ce_9ce_adf_adf_9ce_acd_cef_cef_def_def_ddf_ddf_def_cdf_ace_ace_9bd_9cd_cef_def_cdf_def_def_def_def_def_def_def_def_def_def_def_def_cef_cef_cde_9bc_9cd_cef_bef_9bd_acd_cef_cef_9cd_9cd_ade_9df_9ce_9ce_ace_ace_cdf_def_def_def_def_def_def_def_def_def_def_def_def_def_cef_cdf_9bd_9ce_adf_adf_9ce_9ce_adf_adf_9cf_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8cf_9df_9df_8ce_8ce_9df_9df_8ce_9df_9df_adf_8bd_9cd_def_eef_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_dee_eef_dee_dde_dde_eef_def_eef_eef_eef_def_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eff_cef_8cd_9ce_adf_9df_8ce_8ce_9df_9df_8ce_8df_9df_9df_9ce_9ce_adf_ade_dff_def_def_def_def_def_cef_bef_9cd_9ce_adf_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8df_9df_9df_9ce_ace_dff_eff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eef_eee_eee_eee_eee_eef_eee_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_cef_cef_def_def_cef_bef_9cd_9cf_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce;
				8'b010110100: horiz=6144'h_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_8df_8df_9df_9df_8df_8cf_9ce_adf_acf_ace_ace_bde_cdf_def_eef_eef_eee_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_def_cff_9ce_9de_8ce_8df_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_8df_9df_9df_8ce_9df_9df_adf_cef_cef_cdf_cde_ddf_def_ddf_def_def_cef_cef_cef_cef_cef_cef_bdf_cef_cef_cdf_bdf_cef_cef_cef_cef_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_def_def_def_def_def_def_ddf_ddf_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_eff_fff_def_cee_bde_adf_ace_ace_ace_ace_ace_9ce_9df_9df_8ce_8df_9df_9df_8df_9df_9df_9df_8ce_8df_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8df_9df_9df_8cf_9df_9df_9df_9cf_9cf_9df_9df_8ce_9de_bef_bef_bdf_cef_cef_bdf_cef_bef_adf_9df_9df_9de_aef_bdf_cef_cef_cef_bdf_cef_cdf_def_ddf_def_def_def_cdf_def_def_cef_bdf_bde_ade_cef_bef_acd_ace_bdf_bef_ade_ade_ade_9df_8df_9df_adf_adf_cef_cef_cef_bdf_cef_cef_cef_bdf_cef_cef_cef_bdf_cef_bef_bef_bdf_9ce_9df_9df_9df_9cf_9cf_9df_9df_8cf_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9cf_ade_bde_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eef_eef_def_def_def_def_eef_eef_eef_eef_def_def_eef_eef_eef_def_bef_9ce_ace_adf_adf_9ce_9df_9df_8df_8cf_8df_9df_9ce_ade_ace_bde_bde_def_dee_eef_eef_eee_eef_def_cee_acd_ade_ade_adf_9ce_8df_9df_9df_8ce_9df_9df_9df_8df_8df_9df_9df_8ce_9df_9df_9df_ace_bde_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_def_bdf_bdf_ade_9df_9df_9df_9df_8df_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8ce;
				8'b010110101: horiz=6144'h_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9ef_8ce_8df_9df_9df_8ce_9ce_adf_bdf_def_def_def_eef_def_eef_eef_eef_eef_dee_fff_eff_eff_eff_fff_eff_eff_fff_fff_fff_eff_fff_eff_dff_9cd_9ce_9df_9df_8cf_8cf_9df_9df_8ce_8df_9df_9df_8ce_8df_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_9cf_9ce_adf_bdf_ace_abd_cef_def_def_def_def_bdf_9ce_9ce_adf_adf_9ce_9ce_9df_adf_9ce_9ce_9df_9df_9ce_9cd_cef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eff_fff_eef_eef_def_def_def_def_dee_def_def_cff_9ce_9ce_adf_9df_8ce_8df_9df_9df_8ce_8df_9df_9df_8ce_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8df_9df_9df_8cf_8cf_aef_9df_8cf_8df_9df_9df_8ce_9ce_9df_9df_9ce_9ce_adf_9df_8ce_8df_9df_8df_8ce_9ce_9de_9df_9ce_9ce_ade_bdf_def_ddf_def_cef_acd_ace_cef_cef_acd_acd_cff_bef_9cd_ace_cff_cef_9cd_ace_cef_cef_9ce_9cf_9df_9df_8df_8ce_9df_9df_9ce_9ce_9df_9df_9ce_9ce_9df_9df_9ce_9ce_9de_9df_9ce_8cf_9df_9df_8ce_8cf_9ef_9df_8cf_8df_9df_9df_8ce_9cf_9df_9df_8cf_9cf_9df_9df_8ce_9cf_9df_9df_8cf_8cf_9df_9df_8ce_adf_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_def_def_ddf_ddf_ddf_def_cef_cef_def_cef_bdf_adf_9df_8ce_8df_9ef_9df_9ce_ace_eff_dff_def_def_dee_eef_fff_fff_fff_fff_fff_eff_eff_eff_dff_cef_9df_9df_8ce_9df_9df_9df_8ce_8cf_aef_9df_8ce_8df_9df_9df_8cf_adf_cef_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eee_eee_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_ddf_def_abd_acd_bef_bef_9ce_8ce_9df_9df_8ce_8df_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9df_8cf_8cf_9df;
				8'b010110110: horiz=6144'h_9df_9df_8cf_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_9cf_9cf_9df_8df_8df_8df_9df_9ce_9ce_9cd_ace_cde_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eff_eff_eff_eff_fff_eff_eff_fff_fff_fff_eff_fff_eff_eff_acd_9ce_adf_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_8cf_9df_9df_9df_9cf_9ce_bef_cef_cef_cef_cef_aef_9ce_9cf_9df_9df_8ce_9df_9df_9df_9cf_9df_9df_9df_9ce_9cd_def_def_def_def_def_def_def_def_def_def_def_dee_dee_dee_dee_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eff_fff_eef_eee_eef_def_def_eee_eee_eef_eef_def_acd_acd_bde_adf_8ce_8df_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_8df_8cf_9df_9df_8df_8cf_9df_9df_8df_8df_9df_9df_8cf_9df_9df_8df_8ce_8df_8df_8df_8ce_8df_9df_9df_9df_9df_9df_adf_bef_cef_cef_bef_9ce_9ce_bef_bef_9ce_9ce_bef_bef_9ce_9ce_bef_bef_9ce_9cd_bef_bdf_9ce_9cf_9df_8df_8df_9df_9df_9df_9df_9df_9df_9df_8ce_9df_9df_9df_9df_9df_9df_9df_8cf_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9ce_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_eef_ddf_def_ddf_def_def_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_def_cdf_bef_adf_9df_8df_8df_9df_9df_ade_bcd_eff_def_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_dff_cef_ade_9df_8cf_8ce_9df_9df_9df_8cf_9df_9df_8df_8cf_9df_9df_9ce_ade_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_eef_eff_eff_fff_fff_fff_fff_eff_fff_eff_fff_eef_def_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_def_def_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_def_cdf_bde_ade_ace_bdf_bef_9df_8ce_8de_8df_8df_8cf_9df_9df_9df_8cf_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_9cf_8cf_9df_9df_9df_8cf_9df_9df_9cf_8cf_9df;
				8'b010110111: horiz=6144'h_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8cf_8cf_adf_9df_8cf_8df_9df_9df_9ce_9ce_cef_def_def_eef_eef_eef_edf_eef_def_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_ffe_fff_eff_eff_def_cef_9cf_9df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8cf_8cf_9df_9df_8ce_7cf_9df_8df_8ce_9ce_adf_adf_9ce_8ce_9df_9df_8ce_8cf_9df_9ef_8cf_8cf_9df_9df_8cf_9df_adf_bdf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_dee_eef_dee_eee_dee_dee_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_fff_eff_dff_dff_ade_9df_8ce_8ce_9df_9df_8ce_9df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8ce_9df_9df_9df_8ce_8ce_9df_9df_8ce_9cf_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8cf_8df_9ef_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8ce_9df_9df_9df_9ce_8ce_9ef_9df_8ce_8ce_adf_9df_8ce_9cf_adf_9de_8cd_8ce_adf_9de_9ce_9ce_9df_9df_8ce_8df_9df_9df_8cf_8cf_9df_9df_8ce_8cf_9df_9ef_8cf_8cf_9df_9df_8ce_9df_9df_9df_8cf_8ce_9df_9df_8ce_9df_9df_9df_8ce_8ce_9df_9df_8ce_8df_9df_9df_8ce_8cf_9df_9df_8cf_8df_9df_8df_8ce_9df_adf_bde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_fff_eff_fff_fff_fff_eff_acd_ade_9ce_8ce_9df_9df_8ce_ace_dff_eef_eef_eef_eef_eef_eef_eee_fff_eff_eff_eff_fff_fff_fff_fff_eef_def_9ce_8ce_9df_9df_8ce_8ce_9df_9df_8ce_9df_9df_9df_8ce_9cf_adf_bdf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_fff_fff_fff_eff_dee_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_def_eef_def_eef_eef_eef_eef_eef_eef_ddf_ddf_def_ddf_def_cdf_9cd_9cd_cff_cef_ace_9ce_adf_9df_8ce_8df_9df_9df_8ce_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8cf_9df_9df_9df_8cf_8cf_9df_9df_8cf_9df_9df_9df_8cf;
				8'b010111000: horiz=6144'h_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8ce_9ce_9ce_9df_9df_9cf_9df_8df_9de_ace_bce_def_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_fff_fff_fff_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_dee_dff_9cd_8de_8df_9df_9ce_9cf_adf_9cf_9df_9de_9df_9df_8de_9df_9df_8cf_8cf_9df_9df_9df_9de_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8cf_8cf_9df_9df_9df_9df_8cf_9df_9df_8cf_9cf_9df_9df_9cf_9df_9df_8cf_8cf_9cf_9df_9df_9cf_9df_9df_9cf_9cf_ace_bde_cde_def_eee_eef_eef_eef_eef_eef_eef_eef_def_eef_eff_eff_fff_fff_fff_fff_fff_eee_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_bdd_bef_9cd_8df_9df_8df_8df_8ce_9df_9df_9df_9df_adf_9cf_9ce_9cf_9df_9df_9de_9df_9df_8ce_8ce_9de_9df_9df_9de_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_9cf_9cf_9cf_9df_9df_9cf_8df_9df_8ce_8ce_9df_9df_9df_9cf_9df_9df_8cf_8ce_9de_9de_9df_9de_9df_9df_8cf_8cf_9df_9df_9df_9df_9df_9df_9df_8ce_8df_8df_9df_9df_9df_9df_8cf_8cf_9cf_9df_9df_9cf_9df_9df_8cf_8cf_9df_9df_9df_9de_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8cf_8cf_8df_9df_9df_9ce_9ce_bde_cde_eef_eef_def_def_eef_eef_eef_eef_eef_eee_eee_eee_eff_fff_fff_fff_fff_fff_eee_eff_eef_eef_eef_eef_eef_eef_eef_eef_edf_eef_eef_ddf_def_dde_dde_dde_eef_dee_dee_dee_eff_eff_eff_eff_eff_eff_bdd_bef_8ce_8df_9df_9ce_ade_ccd_eef_eef_eef_eef_eef_eef_eef_eee_fff_eff_fff_fff_fff_fff_fff_fff_eef_def_bcd_ade_adf_9df_9df_9df_9df_9df_8ce_8cf_9df_9df_9df_8df_9df_ade_def_eef_eef_eef_eef_def_def_def_def_def_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_def_def_ddf_def_def_def_eef_eef_eef_eef_eef_eef_ddf_def_bdf_bef_bef_bef_ace_ace_bef_aef_9ce_8df_9df_9df_8ce_9cf_9cf_9df_9df_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8ce_8ce_9df_9df_9df_9df_9df_9df_8ce_8ce_9df_9df_9df_9df;
				8'b010111001: horiz=6144'h_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9de_cef_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_fff_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_dff_ade_9df_9df_9df_9df_9df_8ce_9cf_9df_9df_9df_adf_9df_9df_8ce_9cf_9df_9df_9df_9df_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_8cf_9df_9df_9df_adf_9df_9df_8ce_9cf_9df_9df_9df_9df_9df_9df_8ce_9cf_9df_9df_9df_9df_9df_9df_8cf_9cf_adf_adf_dff_def_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_efe_fff_fff_fff_fff_eff_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_dff_ade_9df_8ce_9ce_adf_9df_9df_adf_9df_adf_9ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9ce_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_8df_9df_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_8cf_9df_9df_9df_9df_9df_9df_8cf_8ce_9ef_9df_9df_9df_9df_9df_8ce_8cf_9df_9df_9df_adf_9df_9df_8cf_9cf_adf_9df_9df_adf_9df_9df_8ce_8df_9df_9df_9df_adf_9df_9df_8ce_9cf_9df_9df_9df_adf_adf_adf_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eff_eff_eff_eff_eff_fff_eff_dff_9de_9df_8ce_ace_dff_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_fff_fff_fff_fff_fff_fff_fff_fff_def_cef_ade_adf_adf_adf_9ce_9ce_adf_9df_9df_9df_9df_9df_8ce_9cd_def_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_def_ddf_def_def_def_ddf_ddf_ddf_def_def_eef_eef_eef_eef_edf_eef_def_ace_9ce_9ce_9ce_adf_acf_adf_9df_9df_9df_8cf_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_8ce_9cf_adf_9df_9df_adf_9df;
				8'b010111010: horiz=6144'h_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9ce_ace_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_dff_ade_9df_9df_adf_adf_8df_8ce_8df_9df_9df_9df_adf_adf_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9df_9df_9df_9df_9df_9df_9df_8ce_9cf_9df_9df_9df_9df_9df_9df_9cf_9df_9df_9df_9df_9df_9df_9df_9cf_9cf_adf_adf_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_eff_fff_fff_fff_fff_eff_eff_bde_ade_9cd_9ce_ade_adf_adf_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9ce_9de_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_adf_9df_9df_8df_9df_9df_9df_9df_adf_adf_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_8df_9df_9df_9df_9df_9df_9df_9df_8cf_8ce_aef_9df_9df_9df_9df_9df_8cf_9df_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9df_9df_9df_9df_adf_9df_9df_9ce_9ce_adf_9df_9df_adf_adf_ace_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_efe_eff_fff_eff_eff_eff_fff_fff_eff_bde_bde_acd_bce_def_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_def_cef_bce_bde_bde_ade_ace_9ce_adf_9df_9df_9df_9df_8df_9de_9cd_def_eef_def_eef_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_eef_eef_eef_def_def_def_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_ddf_def_def_ddf_def_def_ddf_def_def_def_def_def_eef_eef_eef_eef_eef_def_bce_adf_9ce_9bd_adf_adf_9cf_9df_9df_9df_8ce_9cf_adf_9df_9df_adf_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df_9df_9cf_9cf_9df_9df_9df_9df_9df;
				8'b010111011: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_ade_bde_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_fff_eff_dee_dff_ace_ade_9de_adf_ade_adf_adf_9df_9df_9df_9df_adf_9df_adf_adf_9df_adf_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_fff_fff_fff_fff_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_fff_fff_fff_eff_def_def_cef_cef_adf_ace_9df_9df_9df_adf_9cf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_adf_adf_9df_9df_9df_9df_adf_9df_bde_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_dde_eee_eff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_fff_fff_fff_fff_fff_fff_fff_efe_eff_fff_fff_eff_eff_ffe_fff_fff_fff_eff_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_fff_fff_eee_eef_def_def_def_def_fff_eff_dff_cef_ace_ade_9df_adf_9df_9df_9df_ade_def_def_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_def_def_ddf_def_def_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_ddf_eef_eef_eef_eef_def_def_cef_cff_bdf_bdf_cef_cef_adf_9df_aef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b010111100: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_bde_bdf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eff_eff_eff_fff_fff_fff_fff_eff_def_cef_bce_ade_ade_ace_ade_bdf_ade_bdf_ade_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_dff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_efe_fff_fff_fff_fff_fff_eef_eef_def_cdf_bdf_bdf_adf_aef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_ade_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eee_eef_eef_eef_eef_eee_fff_eff_def_def_bdd_bde_ade_adf_9df_9df_adf_ace_def_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_def_def_def_def_def_ddf_ddf_def_def_def_eef_def_eef_eef_eef_eef_eef_eef_eef_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_ddf_def_def_def_def_def_eef_eef_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_ddf_ddf_ddf_def_def_def_def_def_def_def_eef_eef_eef_eef_def_def_cef_bce_bde_def_cdf_bde_bdf_ade_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b010111101: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_dff_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_dee_fff_fff_fff_fff_fff_eff_def_def_def_def_def_def_dff_def_def_def_ace_ade_9de_9df_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_ade_bce_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_eee_eef_eef_eef_def_def_def_cff_ade_ace_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_ade_bde_bcd_eef_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_dee_eef_eef_eef_eef_eef_eef_dee_fff_fff_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_eff_fff_fff_fff_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_eee_eef_eef_dee_eef_eef_eef_eee_fff_eff_fff_eff_def_def_bde_ace_adf_adf_adf_ace_cef_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_def_def_def_def_def_def_def_def_ddf_ddf_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_ddf_ddf_def_def_def_def_def_def_def_def_cef_ade_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b010111110: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_ade_acd_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_eff_eff_eff_eff_eff_def_eef_eef_eef_eef_eef_eff_eee_eef_dde_bdd_bde_ade_ade_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_adf_adf_bde_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_fff_fff_fff_fff_fff_fff_def_eef_eef_eef_eef_def_def_cef_bde_ace_ace_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_adf_bde_bce_bcd_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_eff_eff_eff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_fff_fff_eff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_def_def_bce_ace_bde_adf_adf_ace_cdf_cdf_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_cdf_ace_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b010111111: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_ade_bde_dff_def_eef_eef_eef_eef_def_eef_eef_eee_eee_eef_fff_fff_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_eff_eff_eff_eff_eff_dff_acd_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_adf_bdf_def_eef_eef_eef_eef_eef_eef_eef_eef_edf_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eee_eee_eee_eee_eee_eee_eee_eee_fff_fff_eff_fff_eff_fff_fff_eff_def_eef_eef_eef_eef_eef_dee_def_def_def_cef_cff_ade_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_adf_9df_9df_adf_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_adf_adf_adf_bdf_dff_cef_def_def_ddf_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eee_eee_fff_fff_eff_fff_fff_fff_fff_fff_eee_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_dee_dee_def_def_def_def_def_cdf_bef_9df_9ce_ace_bde_cef_cef_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_def_def_ddf_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_ddf_def_def_def_def_def_def_def_ddf_def_def_def_def_ddf_def_def_ddf_ddf_ddf_ddf_def_cef_cef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000000: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_bdf_cce_def_eef_eef_eef_eef_eef_eef_eee_eee_eee_eef_eef_fff_fff_fff_fff_fff_eff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_fff_fff_fff_fff_fff_fff_fff_def_bdd_bdf_ade_9de_9ef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_cef_def_eff_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_eef_eef_fff_fef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eff_eff_fff_fff_eff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cef_bef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_9df_9df_adf_adf_ade_bdf_bce_bce_bce_bce_adf_adf_9df_9df_9df_9df_9df_adf_acf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_bde_bce_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_eff_eef_eef_eef_def_def_eef_def_eef_def_def_def_def_def_eef_eef_eef_eef_eef_eef_def_def_eef_eef_eef_def_def_def_def_def_cef_cef_cef_cef_cef_cef_aef_adf_9df_9de_adf_bef_cef_cef_cde_def_def_def_ddf_ddf_ddf_ddf_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_eef_ddf_def_cdf_cef_cdf_bdf_cef_def_ddf_edf_edf_ddf_def_def_def_def_def_def_def_def_ddf_def_def_def_def_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bef_bef_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000001: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_bde_dff_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_fff_fff_fff_fff_fff_ffe_efe_fff_fff_fff_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_eff_eff_fff_fff_fff_fff_fff_fff_eff_eff_dff_acd_ade_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_ade_adf_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_ade_bcd_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_fff_fff_fff_eff_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_def_bcd_ade_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_adf_adf_bde_dff_def_def_def_def_cef_adf_ace_adf_adf_adf_adf_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_ade_dff_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_edf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_fff_fff_fff_fff_eee_eef_eef_dee_eef_eef_dde_eef_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_cdf_cef_cef_ade_ace_ade_ade_ade_ace_ace_adf_9df_9df_9df_9de_9de_adf_ace_bce_cef_cdf_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_def_def_def_def_ddf_ddf_def_def_def_ace_ace_bdf_ace_cef_cdf_cdf_ddf_ddf_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_cef_cef_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_ade_adf_adf_adf_aef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000010: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_adf_bde_dff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_efe_eff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eee_fff_fff_fff_eff_fff_fff_fff_fff_fff_eff_eff_dff_bdd_bde_ade_bdf_adf_adf_9df_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_adf_9ce_ade_ace_ace_ace_ace_ace_ace_adf_adf_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_adf_adf_ade_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cde_bde_bde_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_bdf_bde_bde_cde_eef_def_def_def_def_cdf_bce_bce_bce_ace_ace_ace_ace_adf_adf_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_ace_ade_ace_bde_bde_def_eef_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_eff_eef_eef_eef_eef_eef_eef_ddf_def_cdf_cdf_def_ddf_def_def_def_def_cef_cef_cef_cef_def_def_def_ddf_ddf_def_def_def_cef_bef_adf_9ce_adf_9df_9df_9df_adf_9df_adf_9df_9df_9df_9df_adf_adf_bdf_cef_cef_cef_cef_cef_cef_cef_cdf_def_ddf_def_def_def_def_def_def_cef_cef_cef_cdf_def_ddf_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_cef_cdf_cdf_cef_def_cef_cdf_bdf_ade_adf_bdf_cef_cef_cef_cef_cef_cef_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_cdf_cef_cef_cef_cef_cdf_bdf_bef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000011: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_bde_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_eff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_eff_eff_eff_eff_fff_fff_fff_fff_fff_eff_eff_eff_eff_eff_def_def_cef_cef_ade_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_adf_ade_bde_def_def_def_def_def_def_def_cef_ace_adf_adf_9df_9df_adf_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_adf_ade_ace_bde_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_eee_eee_eee_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_dff_cef_ade_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_bdf_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_def_def_cff_ade_ade_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_bce_cef_cef_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_acd_bde_cef_ddf_ddf_def_def_cef_ade_9ce_ade_ade_cef_def_def_def_def_def_def_cef_ade_adf_adf_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bde_cef_cef_def_def_def_cef_cef_cef_ace_ace_ade_bde_cef_cef_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_cef_ace_bde_cef_cef_ace_bde_cef_bef_ade_ade_ade_adf_9df_9ce_ade_ade_cef_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_ddf_def_def_def_cdf_bce_adf_adf_adf_adf_ace_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000100: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9cf_adf_bdf_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_eff_efe_fff_fff_fff_fff_fff_eef_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eff_eff_fff_eef_eef_ddf_cef_bde_adf_adf_adf_9df_9df_9df_9df_9df_adf_bef_ade_bde_bce_def_eef_def_eef_eef_eef_def_cde_bde_bde_ace_adf_9de_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_cef_def_def_def_eef_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_eef_eef_eef_cef_bde_bdf_ade_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_bdf_cef_cef_cef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_cef_bef_ade_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_bce_cdf_cdf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_cef_ade_ade_bef_cef_cef_def_cef_bef_adf_9df_9df_adf_bef_def_def_def_cef_cef_cef_bef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_bde_bdf_cef_cef_cef_cef_cef_cef_bdf_adf_adf_9ce_adf_bef_cef_cef_cef_cef_cef_def_cde_ddf_ddf_ddf_cdf_cdf_def_def_def_def_cef_bde_bde_cef_bdf_bde_bdf_cef_bdf_bdf_bdf_adf_9df_9df_9df_9df_adf_bef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000101: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_ace_bcd_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dde_dee_fff_fff_fff_fff_fff_fff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_def_dff_dff_cef_ade_ade_ade_ade_ade_ade_cef_dff_def_eef_eef_dee_fff_fff_fff_fff_fff_eff_eff_eff_cef_cff_ade_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_ace_bce_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_def_def_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_eff_eff_eff_def_cef_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_ade_ade_ace_acd_bce_def_def_eef_def_def_eef_eef_def_def_def_acd_ace_ade_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_ace_cdf_cdf_cdf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_ddf_ddf_ddf_ddf_ddf_ddf_bdf_ade_9de_9de_9de_adf_ace_adf_adf_adf_aef_9df_9df_9de_9ce_ade_ade_adf_adf_adf_adf_aef_aef_9df_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9ce_adf_adf_ade_ade_ade_adf_adf_adf_9df_adf_9df_9ce_adf_adf_ade_9de_ade_ade_ade_ace_cdf_ddf_ddf_cef_bce_bce_cef_cef_ace_ace_cef_cef_ace_bde_cef_cef_ace_adf_cef_bef_adf_9df_9df_9df_9df_9de_ace_adf_adf_adf_adf_adf_adf_adf_adf_ade_ade_ade_ade_adf_adf_aef_aef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000110: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9ce_ace_bce_bcd_cde_def_eef_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_fff_eff_eff_fff_fff_eff_fff_fff_eee_eef_eef_eef_eef_eef_eef_eef_eff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_cef_bde_ace_ace_ace_ace_bcd_cef_eef_eef_eef_eee_dde_fff_fff_fff_fff_fff_fff_fff_eff_def_cef_ade_9de_adf_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9de_adf_ace_bde_cdf_def_ddf_def_def_def_def_ddf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_eef_ddf_def_ddf_def_def_def_def_ddf_eef_def_eef_def_def_def_def_eef_eef_eef_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_fff_eef_def_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9de_9de_ade_cef_def_def_def_cef_def_def_def_def_bef_ade_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_bef_cef_cef_cdf_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_def_def_ddf_def_def_eef_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_ddf_def_def_def_def_def_def_ddf_eef_def_eef_eef_eef_eef_eef_def_def_def_ddf_def_def_def_def_cef_cdf_bdf_9de_9df_9df_9df_9df_adf_adf_adf_aef_9df_9df_9df_9df_adf_9df_9df_9df_adf_adf_adf_aef_9df_9df_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_adf_adf_cef_cef_cef_cef_bdf_ace_bef_bef_ade_ace_bef_bef_ade_ade_cef_bef_ade_adf_bef_bef_adf_9df_9df_9df_9df_adf_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_aef_aef_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011000111: horiz=6144'h_9df_9df_9df_9df_9df_9df_9df_9df_9de_9de_adf_adf_ace_dff_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_def_dee_dee_dee_eee_fff_fff_dde_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eee_eee_eee_eee_eee_eee_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_def_def_def_eef_eef_eef_eef_eef_eef_def_def_def_def_eef_def_eef_eef_ede_eee_eee_eff_fff_fff_fff_fff_ffe_fff_fff_dee_cff_ade_9de_aef_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9de_adf_cef_cef_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_dde_dde_ddf_ddf_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_eff_fff_fff_fff_fff_fff_eef_def_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9ef_9df_9df_9de_9de_adf_ade_adf_adf_ade_adf_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9ce_adf_ace_bde_def_ddf_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_dde_dde_ddf_ddf_def_ddf_def_ddf_def_def_def_def_def_def_bdf_ace_adf_adf_9df_9df_9df_9df_9df_adf_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_adf_adf_9de_9df_9df_9de_adf_adf_9de_9de_9df_adf_adf_adf_adf_adf_9df_adf_adf_adf_9df_9df_adf_adf_adf_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011001000: horiz=6144'h_9df_adf_adf_9df_9df_9df_9df_adf_adf_adf_ade_bde_bce_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_fff_fff_fff_fff_fff_fff_fff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_fff_fff_fff_eff_eee_def_bcd_bdf_9ce_9df_9df_9df_9df_9df_9df_9df_adf_adf_adf_9df_9df_9df_adf_adf_cdf_def_def_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_ddf_def_cef_def_ddf_def_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_fff_fff_fff_fff_fff_dee_def_bdd_bde_ade_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_bef_cef_bef_cef_cef_cef_cef_cef_cef_cdf_def_def_def_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_dde_def_cdf_bce_bdf_adf_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df;
				8'b011001001: horiz=6144'h_9df_9df_adf_9df_9df_9df_9df_adf_adf_ade_bde_dff_eef_def_eef_fef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_dee_def_eef_eef_eef_eef_eef_eef_eef_def_eef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_fff_eff_def_cef_ace_ade_9de_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_bdf_cef_def_ddf_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_def_def_def_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_fff_fff_fff_fff_fff_eff_fff_eff_dff_cff_ade_9de_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9cf_adf_adf_adf_ade_ade_adf_ade_ade_ace_acd_cef_ddf_def_def_ddf_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_ddf_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_ddf_ddf_ddf_ddf_ddf_cdf_def_cdf_cde_cdf_cef_cef_cef_adf_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df;
				8'b011001010: horiz=6144'h_9df_9df_adf_9df_9df_9df_adf_bdf_bce_bde_bde_eff_eef_eef_eef_eff_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_eff_fff_eff_def_def_def_eef_eef_eef_eef_eef_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_eff_fff_eff_eff_def_def_bde_ace_bde_ade_ace_adf_ade_9df_9df_9df_9df_9df_9df_adf_adf_bdf_cdf_cdf_def_def_def_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_fff_fff_fff_fff_fff_fff_eff_eff_def_cef_bde_ade_ade_bdf_adf_adf_adf_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_adf_adf_adf_9df_9df_9de_9df_9de_9de_bef_cdf_def_def_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_def_def_def_def_def_def_def_def_cef_cef_cef_cef_cef_cef_bef_bef_adf_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_adf_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df_9df_9df_adf_9df_9df_9df_9df_9df;
				8'b011001011: horiz=6144'h_9df_aef_adf_9df_9df_9de_adf_cef_def_eff_def_eef_eef_dee_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_def_def_def_bdf_cdf_bce_bde_def_def_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eee_eef_fff_fff_fff_eff_dee_eee_def_def_def_def_eff_eff_def_dff_bdf_aef_9df_9df_9df_9df_9df_9df_adf_bdf_ade_bce_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_fff_dee_eef_def_def_def_def_eff_eff_dff_cef_ade_adf_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_adf_9df_9df_aef_9df_aef_aef_9de_9ef_adf_9de_9de_bce_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_ddf_def_cdf_cef_cef_ace_ade_ade_ade_bdf_bdf_adf_adf_adf_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_adf_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_adf_aef_adf_9df_9df_9df_9df_9df_adf_aef_adf_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df_9df_aef_aef_9df_9df_9df_9df_9df;
				8'b011001100: horiz=6144'h_9df_adf_aef_adf_adf_ade_ace_def_def_eef_eef_eef_eef_eef_eef_eef_def_def_eef_eef_def_eef_eef_eef_def_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_def_def_def_def_def_cef_bdf_bdf_ade_bde_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_fff_fff_fff_eff_eef_eef_eef_eef_eef_dee_eff_eff_eef_def_cde_bdf_9de_9df_9df_9df_adf_9df_aef_adf_9de_adf_bef_cef_cef_cde_def_def_ddf_ddf_ddf_def_cdf_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cdf_cdf_def_def_ddf_ddf_ddf_def_ddf_ddf_ddf_def_ddf_dde_ddf_def_def_def_def_cde_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_eee_eef_eef_eef_eef_dee_fff_eff_def_def_bce_adf_adf_adf_9df_adf_aef_adf_9df_adf_9df_9de_adf_adf_aef_adf_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_aef_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_bdf_cef_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_ddf_ddf_ddf_ddf_def_cef_cdf_cdf_cef_cef_cde_def_def_ddf_ddf_ddf_def_ddf_ddf_ddf_def_ddf_ddf_ddf_def_def_cef_cef_cef_bef_bef_adf_9df_adf_adf_adf_aef_adf_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_9df_adf_aef_adf_adf_adf_9df_adf_adf_aef_adf_adf_adf_9de_adf_adf_adf_aef_adf_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef_adf_adf_aef_9df_adf_9df_9df_aef;
				8'b011001101: horiz=6144'h_aef_9df_adf_aef_adf_adf_ade_cef_ddf_ddf_def_dde_ddf_ddf_ddf_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_ddf_ddf_ddf_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_ddf_ddf_ddf_ddf_ddf_cdf_bde_ade_ade_ace_bdf_bdf_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eee_eef_eef_eef_eef_eef_eef_dee_fff_fff_fff_fff_def_def_bdf_bef_adf_adf_bdf_aef_9df_9df_aef_aef_9de_ade_adf_bde_cef_def_def_ddf_cdf_cef_bdf_adf_ace_ade_adf_adf_ace_ade_adf_adf_9de_ade_bdf_bdf_cdf_def_def_ddf_cdf_def_def_ddf_cdf_def_def_cef_cdf_def_def_cef_bce_bce_dff_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eef_eef_eee_eef_eef_def_eef_eef_eef_eee_fff_eff_fff_eff_def_cef_ade_ade_bef_bef_ade_adf_aef_aef_adf_adf_aef_aef_9de_9df_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_aef_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_aef_9ce_adf_bef_aef_9df_9df_aef_adf_9ce_adf_bef_aef_9df_adf_bef_bdf_ace_bce_def_ddf_ddf_ddf_def_ddf_ddf_def_def_def_def_def_def_ddf_def_cef_bdf_bdf_ace_adf_bdf_cde_cdf_def_def_cdf_cdf_def_def_cdf_cdf_def_ddf_ddf_cdf_def_def_cef_acd_adf_adf_adf_9df_9df_aef_aef_9df_adf_aef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_adf_9df_adf_aef_bef_ade_ade_bef_bdf_adf_adf_aef_aef_9df_adf_aef_adf_9de_adf_aef_aef_9de_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef_adf_9ce_adf_bef_aef_9df_adf_aef;
				8'b011001110: horiz=6144'h_aef_adf_adf_adf_adf_adf_adf_bdf_cef_cef_cef_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_eef_def_eef_eef_eef_eef_eef_def_def_eef_eef_eef_eef_eef_ddf_def_def_def_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_ddf_ddf_ddf_def_def_cef_bde_bef_ade_ade_ade_bdf_cef_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_fff_fff_fff_eff_def_def_cdf_cdf_bde_ade_adf_adf_adf_9de_aef_9df_9df_adf_adf_bdf_cef_cef_cef_cef_cef_cef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_9df_adf_adf_bdf_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bef_ade_ade_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eee_fff_fff_fff_fff_eef_def_bde_bde_cef_bdf_ade_ade_adf_adf_adf_adf_adf_adf_adf_adf_aef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_aef_ade_bde_def_def_ddf_def_def_ddf_ddf_def_cef_cef_cef_cef_def_cef_cef_bef_adf_adf_9df_adf_adf_bdf_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bef_ade_adf_adf_adf_adf_adf_adf_aef_adf_9df_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_9df_adf_adf_bdf_bdf_ace_cef_cef_bde_adf_adf_adf_adf_adf_aef_adf_9df_adf_aef_adf_adf_adf_aef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf_adf_9df_adf_bef_adf_adf_adf_adf;
				8'b011001111: horiz=6144'h_ade_aef_adf_adf_9df_aef_bdf_ace_ace_bdf_bdf_cef_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_def_def_def_def_def_def_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_ddf_ddf_def_def_cef_cef_bdf_bdf_9ce_ade_bdf_cdf_def_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eee_eef_eef_eef_eef_eef_eef_eef_def_bdf_ade_bdf_bef_adf_9df_adf_aef_adf_adf_ade_adf_bdf_ace_ace_adf_bdf_adf_adf_aef_aef_9df_adf_aef_aef_9df_adf_aef_adf_adf_9de_adf_adf_9de_ace_adf_adf_ace_ace_adf_adf_ace_ace_adf_bdf_ace_adf_adf_aef_ace_bce_def_eef_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dee_eee_eee_eef_eef_eef_eef_def_def_def_cef_bef_adf_ace_ade_bdf_bef_9ce_ade_aef_aef_9ce_adf_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_ade_adf_aef_9df_9df_aef_aef_9df_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_adf_adf_adf_aef_aef_9de_ade_aef_aef_9df_adf_aef_adf_9cf_9df_aef_aef_9df_9df_aef_aef_9df_9df_bef_bef_def_def_def_def_def_ddf_def_def_cef_cef_bde_cde_def_cdf_bde_adf_9df_9df_aef_aef_9df_9de_adf_adf_ade_9ce_adf_adf_ace_9ce_adf_adf_ace_ace_adf_adf_9de_9df_aef_adf_9df_9df_adf_aef_9de_adf_aef_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_adf_adf_adf_aef_aef_9de_adf_adf_adf_adf_adf_aef_aef_9de_9df_aef_aef_9df_9df_adf_aef_adf_bde_dff_def_dff_dff_def_bdf_ace_adf_bef_adf_adf_adf_aef_adf_adf_9de_aef_aef_9ce_adf_aef_adf_9ce_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de_adf_adf_aef_9df_9df_aef_aef_9de;
				8'b011010000: horiz=6144'h_adf_aef_adf_9de_adf_aef_adf_9cf_adf_adf_bdf_cef_cef_cef_cef_cdf_cef_cef_cef_bef_cef_def_def_dde_ddf_ddf_ddf_def_def_def_def_def_def_def_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_def_ddf_ddf_def_def_cef_cef_cef_def_def_ddf_cde_bdf_9ce_adf_ade_bde_def_eef_eef_eef_eef_eef_eef_def_def_eef_eef_eef_def_def_def_eef_ddf_eef_eef_def_def_eef_def_def_eef_eef_eef_eef_eef_def_def_def_cce_cde_cdf_bdf_bde_adf_bdf_bdf_acf_adf_bdf_adf_9ce_adf_aef_aef_9de_adf_aef_adf_9df_adf_adf_aef_9df_adf_aef_adf_9df_adf_aef_aef_9de_adf_aef_adf_9df_adf_aef_aef_9de_adf_aef_adf_9df_adf_aef_adf_9ce_cde_def_def_eef_eef_eef_eef_def_def_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_eef_def_eef_def_def_ddf_cee_cde_cde_bde_bde_bdf_cef_bdf_adf_bef_adf_adf_adf_adf_bdf_ace_adf_adf_aef_9de_adf_aef_aef_9de_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_aef_adf_9de_adf_aef_aef_9de_adf_adf_bdf_bef_cef_bef_cef_cef_cef_cef_cef_cef_cef_bdf_bdf_cef_bef_bef_aef_adf_adf_aef_aef_9de_adf_aef_adf_9df_adf_aef_adf_9df_adf_aef_adf_9df_adf_aef_aef_9de_adf_aef_adf_9de_adf_adf_adf_adf_adf_aef_adf_9df_adf_aef_aef_9de_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_aef_aef_adf_9de_adf_bef_adf_ade_adf_bef_adf_9ce_ade_adf_bdf_ade_adf_aef_adf_9de_adf_adf_aef_9de_adf_aef_adf_adf_adf_aef_adf_9cf_adf_adf_aef_9de_aef_aef_ade_bdf_cde_def_def_def_def_def_def_cce_cde_cdf_bde_bde_bdf_adf_bdf_acf_adf_bdf_bdf_ace_adf_bdf_adf_9de_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce_adf_bef_adf_9de_adf_aef_adf_9ce;
				8'b011010001: horiz=6144'h_aef_9de_9de_bef_adf_9de_adf_aef_aef_9ce_adf_bef_bdf_ace_bdf_bdf_bdf_ace_adf_bdf_bdf_cef_def_ddf_ddf_ddf_ddf_def_def_def_def_def_ddf_ddf_ddf_def_def_ddf_ddf_def_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_def_cef_cef_cdf_def_def_def_cef_cef_adf_adf_9de_ade_cef_ddf_def_def_ddf_ddf_def_def_def_def_ddf_def_def_def_ddf_def_ddf_ddf_ddf_ddf_def_def_def_def_eef_eef_eef_eef_eef_eef_def_eef_def_eef_eef_def_cef_cef_ade_ade_bef_aef_9df_9df_adf_aef_adf_9df_aef_aef_9df_9df_aef_adf_9ce_adf_bef_aef_9df_9df_bef_aef_9df_9df_aef_aef_9df_9df_aef_aef_adf_9df_adf_bef_9df_9df_aef_aef_adf_adf_adf_bde_cdf_def_def_ddf_ddf_def_ddf_ddf_ddf_def_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_dde_dde_ddf_ddf_ddf_ddf_ddf_ddf_def_eef_eef_eef_def_def_def_cef_cef_bdf_aef_9ce_adf_bef_bef_adf_adf_adf_aef_9df_adf_aef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_aef_9df_9de_aef_aef_adf_adf_adf_aef_9ce_ace_bdf_bdf_ace_adf_adf_bdf_ace_adf_bdf_bdf_ade_ade_bdf_adf_adf_adf_adf_aef_adf_9df_aef_aef_9df_9df_aef_aef_9df_9df_aef_aef_9df_9df_aef_aef_9df_9df_aef_aef_9df_9de_aef_aef_9ce_adf_bef_aef_9df_9df_aef_aef_adf_9df_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_aef_9df_9de_bef_bef_ade_ade_bef_aef_9de_adf_aef_bef_adf_adf_aef_adf_9ce_adf_bef_aef_ade_adf_aef_aef_9de_9de_aef_aef_adf_adf_adf_adf_adf_adf_aef_aef_adf_bde_dff_eef_def_eef_eef_eef_def_eef_eef_def_eef_def_cef_cef_ade_ade_bef_aef_9de_adf_bef_bef_adf_adf_adf_aef_9df_9de_aef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf_bef_adf_9de_bef_aef_adf_adf_adf;
				8'b011010010: horiz=6144'h_aef_adf_9df_adf_adf_adf_9df_aef_aef_9df_9df_aef_adf_adf_adf_adf_adf_adf_adf_adf_bdf_cef_cef_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_def_def_def_ddf_ddf_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_def_cdf_cef_cef_cef_cef_cdf_cef_bef_adf_aef_adf_ade_cef_cdf_cef_cef_def_def_def_def_def_def_cef_cef_cdf_cdf_def_def_def_ddf_ddf_def_def_ddf_def_eef_eef_eef_eef_eef_eef_eef_def_def_def_eef_eef_def_def_def_ade_9de_aef_9ef_9ef_9de_aef_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_adf_bef_adf_adf_9df_aef_aef_adf_9df_aef_aef_adf_9df_adf_adf_adf_9df_adf_adf_adf_9df_aef_adf_adf_9de_adf_bdf_cdf_cef_cdf_cdf_def_def_def_def_ddf_def_cdf_cef_cef_ddf_ddf_def_def_def_def_def_ddf_ddf_def_eef_eef_def_def_def_def_def_eef_eef_eef_eef_eef_def_def_def_bef_bef_ade_adf_aef_adf_adf_9df_aef_aef_adf_9de_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_9df_9ce_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_9df_adf_adf_adf_9df_adf_9de_aef_adf_9de_aef_aef_adf_9df_adf_adf_adf_9df_adf_aef_adf_9df_adf_aef_adf_9df_aef_adf_adf_9df_adf_adf_adf_adf_bef_adf_adf_9df_adf_adf_adf_9df_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_aef_adf_9df_adf_9ef_9df_9df_aef_adf_adf_9de_adf_adf_adf_adf_bef_adf_adf_adf_adf_aef_aef_9de_adf_aef_adf_9de_aef_adf_adf_ade_cef_bdf_bde_bde_def_eef_eef_eef_eef_eef_eef_eef_ddf_eef_eef_def_def_def_ade_9de_aef_9ef_9df_9df_aef_adf_adf_ade_adf_adf_adf_9df_aef_aef_adf_9de_aef_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf_adf_adf_9df_adf_adf_adf_9de_adf;
				8'b011010011: horiz=6144'h_9de_aef_aef_9ce_adf_aef_adf_9df_9df_aef_aef_9de_9df_aef_aef_9df_adf_aef_aef_9df_ade_bdf_cdf_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_def_ddf_ddf_ddf_ddf_ddf_def_def_def_ddf_cdf_cdf_ddf_def_def_def_ddf_def_def_def_def_def_def_def_def_def_def_ddf_ddf_ddf_def_def_def_cef_def_cef_ace_ace_ade_bdf_ace_ace_bdf_adf_9df_9df_adf_adf_9ce_ade_bdf_bdf_cef_cef_def_def_def_cef_bdf_bdf_ace_ace_cef_cef_cdf_def_def_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dff_cff_ade_adf_bef_adf_9ce_ade_adf_aef_adf_adf_bef_aef_9ce_adf_adf_adf_9df_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_adf_aef_aef_9ce_9df_adf_aef_adf_ace_bdf_bdf_ace_bce_cef_cef_cef_ddf_def_cef_ace_ade_bdf_cdf_def_def_def_def_def_def_ddf_ddf_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eff_def_cff_bdf_bdf_ade_ade_adf_aef_9df_adf_aef_adf_9df_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_adf_bef_aef_9ce_9df_adf_aef_adf_9df_adf_adf_9ce_9df_aef_aef_9de_9df_aef_aef_9df_9df_adf_aef_9df_adf_aef_aef_9de_9df_adf_aef_9df_9df_aef_aef_9ce_9de_adf_aef_9df_9df_aef_aef_9ce_9df_adf_aef_adf_adf_bef_aef_9ce_9df_adf_aef_9de_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_adf_bef_aef_9ce_9de_aef_aef_9ce_9df_aef_aef_9ce_adf_bdf_bdf_adf_adf_bef_adf_9ce_adf_adf_adf_9df_9ce_adf_aef_9df_9df_adf_aef_9df_adf_bef_cdf_def_def_dff_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_dff_cff_ade_9df_aef_adf_9de_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf_9df_aef_aef_9ce_9df_adf_aef_adf;
				8'b011010100: horiz=6144'h_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_aef_9de_adf_aef_adf_9df_adf_adf_bdf_cdf_cdf_def_def_ddf_ddf_ddf_ddf_def_ddf_ddf_def_ddf_ddf_def_def_ddf_def_cdf_cdf_cef_def_def_def_def_ddf_ddf_def_ddf_def_def_def_def_ddf_def_def_ddf_ddf_def_def_cef_cef_cef_bdf_ade_ade_bef_adf_9ce_adf_bef_adf_9df_9df_aef_aef_9ce_ade_adf_bef_bdf_cef_cdf_cef_cef_bef_bdf_adf_ace_adf_bef_cef_cef_cef_cef_cdf_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_edf_eef_eef_def_bde_bde_bdf_bdf_ade_adf_bef_aef_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_bef_adf_9ce_adf_aef_adf_ade_bdf_bef_cef_cef_cdf_cef_cef_adf_adf_adf_bef_cdf_cef_cdf_cef_cdf_cdf_def_def_eef_def_eef_eef_def_eef_eef_eef_eef_def_eef_eef_eef_eef_eef_eef_eef_cdf_cdf_cdf_bde_bdf_bef_adf_adf_adf_adf_aef_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_9df_aef_aef_9de_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_adf_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_9df_aef_adf_adf_adf_adf_bef_ade_bdf_bdf_cdf_bdf_adf_adf_bdf_adf_adf_aef_adf_9de_adf_bef_adf_9df_9df_aef_aef_9de_adf_bef_bdf_def_def_def_eef_eef_eef_eef_eef_eef_eef_eef_eef_eef_def_eef_eef_edf_eef_eef_def_bde_bdf_bdf_bdf_ade_adf_aef_aef_9de_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce_adf_aef_adf_9df_adf_aef_aef_9ce;
				8'b011010101: horiz=6144'h_aef_9df_9df_bef_aef_adf_adf_aef_bef_9cf_adf_bef_bef_adf_adf_aef_aef_9df_9df_aef_aef_9ce_ade_bdf_cdf_def_def_ddf_ddf_ddf_ddf_def_def_def_def_ddf_def_def_def_cef_def_bce_ace_bdf_bdf_ace_bce_def_ddf_cdf_def_def_def_def_def_def_cef_cef_def_cdf_def_cef_cef_bdf_bef_ade_ace_bef_bef_adf_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9ce_ade_adf_bdf_ace_ade_bdf_adf_9df_adf_adf_aef_ace_ade_bdf_bef_ace_bde_def_cef_def_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_ddf_cde_dde_def_ddf_ddf_ddf_ddf_ddf_ddf_def_cef_bdf_bef_adf_9df_aef_aef_9df_9df_bef_aef_adf_adf_aef_aef_9df_9df_bef_aef_adf_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_bef_adf_adf_aef_aef_9df_9df_bef_aef_ace_ade_bdf_bdf_ade_adf_aef_aef_9de_adf_bdf_bdf_ace_bde_bdf_bdf_cef_cdf_ddf_def_ddf_def_dde_ddf_ddf_def_def_cef_def_def_def_ddf_ddf_ddf_ddf_cef_cdf_cef_cef_cef_adf_ace_bef_aef_9df_adf_aef_aef_adf_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_adf_adf_aef_aef_9df_9df_bef_aef_9df_9df_aef_aef_9df_adf_bef_bef_adf_adf_adf_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_adf_adf_aef_aef_9df_9df_bef_aef_adf_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9de_adf_bef_adf_ace_bde_def_def_def_eef_def_cef_ade_ace_bdf_adf_adf_ade_adf_aef_adf_9de_aef_aef_9df_9df_aef_aef_ade_ace_def_ddf_def_ddf_dde_ddf_ddf_ddf_def_def_ddf_ddf_ddf_dde_ddf_def_ddf_ddf_ddf_ddf_def_ddf_def_cef_bdf_bef_adf_9df_aef_aef_9df_9df_bef_aef_9df_9df_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef_aef_9df_9df_bef_aef_9df_adf_aef;
				8'b011010110: horiz=6144'h_adf_adf_adf_aef_adf_adf_9de_aef_adf_adf_adf_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_9df_9ce_bdf_bde_def_def_ddf_ddf_ddf_def_def_ddf_def_def_cdf_cdf_def_cef_cdf_cef_bdf_ace_bef_adf_adf_ace_bef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_cef_bef_adf_adf_adf_9df_adf_adf_adf_9df_aef_adf_adf_9df_aef_adf_adf_9df_aef_aef_9de_9de_adf_adf_adf_adf_adf_adf_9df_adf_adf_adf_adf_adf_bef_adf_adf_ade_cef_cef_cef_cdf_def_def_def_def_def_def_def_def_def_def_def_def_cdf_cef_cef_def_cef_cdf_cef_cef_adf_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_9df_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_bdf_adf_aef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_cef_cef_cef_cdf_def_def_def_ddf_def_def_def_def_def_def_def_def_cef_cef_cef_cef_cef_cef_bef_bef_bdf_adf_bdf_adf_adf_9df_adf_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_adf_bdf_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_9df_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_9df_aef_aef_adf_ade_cef_bdf_ace_bce_eef_eef_eef_eef_eef_cef_bde_acd_bde_bdf_bde_bdf_bdf_bef_adf_adf_adf_adf_adf_9df_aef_aef_adf_ace_cef_cdf_cef_cef_def_def_def_def_def_def_def_def_def_ddf_def_def_cdf_cef_cef_def_def_cdf_cef_cef_adf_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef_adf_adf_adf_aef_adf_adf_9df_aef;
				8'b011010111: horiz=6144'h_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_adf_aef_aef_9ce_9df_aef_adf_9ce_ade_cef_cef_ddf_ddf_ddf_def_def_def_def_cef_bcd_bce_def_cdf_ace_ace_cef_bef_9df_9df_aef_aef_9de_ace_adf_adf_ace_ade_adf_ade_ace_ade_bde_bde_ace_ace_bdf_adf_9de_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_aef_adf_9de_adf_aef_adf_9de_adf_aef_adf_9de_9de_adf_aef_9df_9df_aef_adf_9df_9df_aef_aef_ace_ace_bdf_bde_def_def_def_def_def_def_def_def_def_ddf_def_cef_ace_ade_bef_bdf_ade_adf_adf_adf_9de_adf_aef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_aef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_ade_aef_aef_9ce_9df_aef_adf_9cf_9df_aef_aef_adf_adf_aef_adf_9df_9df_aef_aef_9de_9de_adf_ade_ace_bce_def_cdf_ddf_def_def_def_def_ddf_def_def_def_cef_bdf_adf_9ce_ade_bef_adf_ade_ade_bef_adf_9ce_adf_adf_adf_9df_adf_bef_adf_9ce_adf_aef_aef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_adf_bdf_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_aef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_bef_adf_9ce_9df_aef_aef_9ce_adf_aef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_aef_9ce_9de_bef_bdf_dff_cef_def_def_dde_eee_eee_eef_eef_eef_def_def_def_eef_eff_def_def_cff_bdf_adf_9ce_adf_bef_adf_9ce_9df_aef_bdf_ace_ade_bdf_bdf_def_def_def_def_def_def_def_def_def_ddf_def_cef_ace_adf_bef_bdf_adf_ade_adf_adf_9ce_adf_bef_adf_9ce_adf_aef_aef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce_adf_aef_bef_9ce_adf_bef_adf_9ce;
				8'b011011000: horiz=6144'h_adf_aef_adf_9de_adf_aef_adf_adf_adf_aef_adf_9de_adf_aef_adf_adf_adf_bef_adf_ade_adf_bef_adf_adf_adf_bef_bef_cef_cef_cef_cdf_def_cef_cef_bdf_bde_bdf_cef_cef_bdf_bdf_cef_bdf_ade_bdf_bdf_adf_ade_adf_bef_adf_9ce_adf_aef_adf_adf_adf_aef_adf_9de_adf_aef_adf_adf_adf_bdf_adf_ace_adf_bef_adf_adf_adf_aef_adf_9de_adf_aef_adf_adf_adf_bef_adf_ade_adf_aef_adf_adf_adf_bef_adf_9ce_adf_aef_adf_adf_adf_aef_adf_9de_ade_adf_bef_cef_cef_bef_cef_cef_cef_cef_cef_cef_cef_cef_bef_adf_adf_aef_aef_9de_adf_aef_adf_9de_adf_aef_aef_9de_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_adf_adf_aef_adf_9de_adf_aef_adf_ade_adf_bef_adf_9ce_adf_aef_adf_adf_adf_aef_adf_9ce_adf_bef_bdf_adf_bdf_cef_cef_cef_cef_cef_cef_cef_cef_bef_bef_bef_bef_bef_adf_9de_adf_aef_adf_adf_adf_bef_bdf_adf_adf_bef_ade_ade_adf_aef_adf_adf_adf_aef_adf_9de_adf_aef_aef_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_bef_bef_cef_cef_cef_cef_def_def_def_def_def_eef_eef_eef_eef_eef_def_def_cef_cff_adf_adf_9ce_adf_aef_adf_adf_adf_aef_adf_9de_ade_adf_bef_bef_cef_bef_cef_cef_cef_cef_cef_cef_cef_cef_bef_adf_adf_aef_aef_9de_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_aef_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade_adf_aef_adf_9de_adf_aef_adf_ade;
				8'b011011001: horiz=6144'h_bef_ade_adf_bef_adf_bef_aef_adf_bef_ade_adf_bef_adf_bef_aef_adf_bef_ade_adf_bef_adf_bef_bef_adf_aef_9de_ade_bdf_bdf_bdf_cdf_cef_cef_ace_bde_cef_cef_ade_bdf_cef_cef_ace_ade_cef_cef_bef_adf_adf_bef_adf_adf_bef_adf_aef_aef_adf_aef_ade_adf_bef_adf_aef_aef_adf_bef_ade_adf_bef_adf_bef_bef_adf_bef_adf_adf_bef_adf_bef_aef_adf_bef_adf_adf_aef_adf_bef_aef_adf_bef_adf_adf_bef_adf_bef_aef_adf_aef_9de_ade_bef_adf_bdf_bdf_bdf_bdf_ace_ade_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bef_adf_aef_aef_adf_aef_9de_ade_bef_adf_aef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_adf_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_adf_adf_bef_adf_aef_aef_adf_aef_9df_9df_bef_adf_bef_bdf_adf_bef_ade_ade_bdf_bdf_bdf_bdf_bdf_bdf_ace_ade_adf_adf_adf_adf_aef_aef_9de_adf_bef_adf_bef_bdf_adf_bef_adf_adf_aef_adf_bef_aef_adf_aef_ade_ade_bef_adf_aef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_aef_9de_ade_bef_bef_adf_bdf_adf_bdf_ace_bde_def_def_def_def_def_def_def_def_def_def_bde_bde_cef_adf_adf_9ce_bef_adf_bef_aef_adf_aef_9df_adf_bef_adf_adf_bdf_adf_bdf_ace_ade_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bef_adf_aef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_aef_ade_ade_bef_adf_aef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf_bef_ade_ade_bef_adf_bef_aef_adf;
				8'b011011010: horiz=6144'h_aef_adf_ade_bef_adf_adf_aef_adf_adf_adf_ade_bef_adf_adf_aef_adf_bdf_adf_ade_bef_adf_adf_bdf_adf_adf_adf_adf_bef_bdf_bdf_bdf_cef_bef_adf_adf_bef_bef_adf_bdf_cef_cef_bde_ade_cef_cef_bef_bdf_bdf_aef_adf_9de_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_adf_adf_ade_bef_adf_adf_bdf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_aef_adf_9ce_bef_adf_adf_adf_adf_aef_adf_ade_bef_bdf_bdf_bdf_adf_bdf_ade_adf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_9de_bef_adf_adf_aef_adf_aef_adf_9de_bef_adf_adf_bdf_adf_adf_ade_ade_bef_adf_adf_adf_adf_adf_ade_adf_adf_bdf_adf_bdf_bef_adf_adf_adf_aef_adf_adf_bdf_adf_adf_adf_adf_adf_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_bdf_adf_bdf_bdf_bde_bde_cef_def_def_def_def_def_def_cef_cef_cef_bef_adf_bef_adf_adf_adf_aef_adf_adf_adf_adf_aef_adf_9de_bef_aef_bef_bdf_adf_bdf_ade_adf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf_aef_adf_ade_bef_adf_adf_aef_adf;
				8'b011011011: horiz=6144'h_bef_aef_adf_adf_adf_adf_aef_adf_aef_aef_adf_adf_adf_adf_aef_adf_bef_bef_adf_adf_adf_adf_bef_adf_bef_bef_adf_bef_adf_bef_bdf_bdf_bef_bef_adf_adf_bdf_bdf_bdf_bef_bdf_bef_adf_adf_bdf_bef_adf_bdf_bef_bef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_bdf_adf_adf_adf_adf_bef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_bef_adf_adf_adf_adf_aef_adf_bef_bef_adf_adf_adf_adf_aef_adf_bef_bef_adf_adf_adf_adf_bdf_aef_bdf_bef_bef_bdf_adf_adf_adf_adf_bef_bef_bef_bdf_adf_adf_bef_adf_bef_bef_adf_adf_adf_adf_bef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_bef_adf_adf_adf_adf_aef_adf_aef_bef_adf_adf_adf_adf_bdf_adf_aef_aef_adf_bef_adf_adf_adf_adf_aef_aef_bef_bdf_bef_bdf_bdf_adf_aef_aef_adf_aef_adf_adf_bdf_adf_bef_bef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_bef_adf_adf_bef_bef_bdf_aef_bef_bef_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_aef_aef_bef_bef_adf_adf_adf_adf_aef_adf_aef_aef_adf_adf_adf_adf_bdf_bef_bdf_bef_bef_bdf_adf_adf_adf_adf_bef_bef_bef_bdf_adf_adf_bef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf_bef_aef_adf_adf_adf_adf_aef_adf;
				8'b011011100: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_aef_aef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_adf_adf_adf_adf_aef_adf_adf_adf_adf_adf_adf_adf_adf_aef_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_aef_aef_adf_adf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_adf_adf_adf_adf_aef_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_aef_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011011101: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_aef_adf_adf_adf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011011110: horiz=6144'h_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf;
				8'b011011111: horiz=6144'h_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_adf_adf_adf_adf_aef_aef_aef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_aef_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_aef_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_aef_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_adf_aef_adf_adf_bdf_bdf_adf_adf_aef_aef_aef_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_aef_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_adf_adf_adf_adf_adf_adf_adf_adf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf_bdf;
				8'b011100000: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100001: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100010: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100011: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100100: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100101: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100110: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011100111: horiz=6144'h_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011101000: horiz=6144'h_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011101001: horiz=6144'h_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011101010: horiz=6144'h_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_adf_adf_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bdf_adf_adf_bdf_bef_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011101011: horiz=6144'h_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bef_adf_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf_adf_bef_bef_bdf_bdf_bef_bef_bef_adf_adf_adf_adf_adf_adf_adf_adf;
				8'b011101100: horiz=6144'h_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_adf_adf_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef_bdf_bef_bef_adf_bdf_bef_bef_bdf_bdf_adf_ade_bef_bdf_adf_ade_bef;
				8'b011101101: horiz=6144'h_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_ade_bef_bef_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef_bef_bef_adf_bef_bef_bef_bdf_bdf_bef_adf_bdf_cef_bef_adf_bdf_cef;
				8'b011101110: horiz=6144'h_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_bef_bef_bef_adf_bef_adf_bef_bef_bef_adf_bef_bef;
				8'b011101111: horiz=6144'h_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_adf_bef_bef_bef_bdf_bef_bef_adf_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf_bdf_bdf_bef_bef_bdf_bdf_bef_bef_adf_bef_bef_adf_adf_bef_bef_adf;
				8'b011110000: horiz=6144'h_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf_bef_bef_bef_bef_bdf_bef_bef_adf;
				8'b011110001: horiz=6144'h_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef;
				8'b011110010: horiz=6144'h_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef_bef_bef_bdf_bef_bef_bef_adf_bef;
				8'b011110011: horiz=6144'h_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef_ade_bef_bef_bdf_adf_bef_bef_bef;
				8'b011110100: horiz=6144'h_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade_bdf_bef_bef_adf_bef_bef_bef_ade;
				8'b011110101: horiz=6144'h_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef;
				8'b011110110: horiz=6144'h_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef_bef_bef_adf_bef_bef_bef_ade_bef;
				8'b011110111: horiz=6144'h_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade_adf_bef_bef_bef_bef_bef_bef_ade;
				8'b011111000: horiz=6144'h_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef_bdf_bef_bef_ade_bef_bef_bef_bef;
				8'b011111001: horiz=6144'h_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef_bef_bef_bde_bef_bef_bef_bef_bef;
				8'b011111010: horiz=6144'h_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef_cef_bef_bde_cef_bef_bef_bef_bef;
				8'b011111011: horiz=6144'h_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef_bef_cef_bef_bef_bef_bef_bef_bef;
				8'b011111100: horiz=6144'h_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef;
				8'b011111101: horiz=6144'h_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef;
				8'b011111110: horiz=6144'h_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef;
				8'b011111111: horiz=6144'h_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef_bef;



                
                default: horiz = 480'h_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00_F00;
            endcase
        end
        else begin
            horiz = 480'h_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0_FF0;
        end
    end
    
endmodule

